module FIR_LPF
(
    input                   clk     ,
    input                   rst     ,
    input                   pls20k  ,
    input   signed [11:0]   din     ,

    output  signed [11:0]   dout
);

    
endmodule 