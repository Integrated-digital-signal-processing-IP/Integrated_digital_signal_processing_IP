module usin_rom
(
input	wire			clka	,
input	wire			rsta 	,
input	wire	[11:0]	addra	,
output	reg 	[11:0]	douta
);
		
always@ ( posedge rsta, posedge clka )
begin
	if ( rsta == 1 )
		douta <= 0;
	else
		case ( addra )
		12'h000 : douta <= 12'h800 ;
		12'h001 : douta <= 12'h803 ;
		12'h002 : douta <= 12'h806 ;
		12'h003 : douta <= 12'h809 ;
		12'h004 : douta <= 12'h80C ;
		12'h005 : douta <= 12'h80F ;
		12'h006 : douta <= 12'h812 ;
		12'h007 : douta <= 12'h815 ;
		12'h008 : douta <= 12'h819 ;
		12'h009 : douta <= 12'h81C ;
		12'h00A : douta <= 12'h81F ;
		12'h00B : douta <= 12'h822 ;
		12'h00C : douta <= 12'h825 ;
		12'h00D : douta <= 12'h828 ;
		12'h00E : douta <= 12'h82B ;
		12'h00F : douta <= 12'h82F ;
		12'h010 : douta <= 12'h832 ;
		12'h011 : douta <= 12'h835 ;
		12'h012 : douta <= 12'h838 ;
		12'h013 : douta <= 12'h83B ;
		12'h014 : douta <= 12'h83E ;
		12'h015 : douta <= 12'h841 ;
		12'h016 : douta <= 12'h845 ;
		12'h017 : douta <= 12'h848 ;
		12'h018 : douta <= 12'h84B ;
		12'h019 : douta <= 12'h84E ;
		12'h01A : douta <= 12'h851 ;
		12'h01B : douta <= 12'h854 ;
		12'h01C : douta <= 12'h857 ;
		12'h01D : douta <= 12'h85B ;
		12'h01E : douta <= 12'h85E ;
		12'h01F : douta <= 12'h861 ;
		12'h020 : douta <= 12'h864 ;
		12'h021 : douta <= 12'h867 ;
		12'h022 : douta <= 12'h86A ;
		12'h023 : douta <= 12'h86D ;
		12'h024 : douta <= 12'h870 ;
		12'h025 : douta <= 12'h874 ;
		12'h026 : douta <= 12'h877 ;
		12'h027 : douta <= 12'h87A ;
		12'h028 : douta <= 12'h87D ;
		12'h029 : douta <= 12'h880 ;
		12'h02A : douta <= 12'h883 ;
		12'h02B : douta <= 12'h886 ;
		12'h02C : douta <= 12'h88A ;
		12'h02D : douta <= 12'h88D ;
		12'h02E : douta <= 12'h890 ;
		12'h02F : douta <= 12'h893 ;
		12'h030 : douta <= 12'h896 ;
		12'h031 : douta <= 12'h899 ;
		12'h032 : douta <= 12'h89C ;
		12'h033 : douta <= 12'h89F ;
		12'h034 : douta <= 12'h8A3 ;
		12'h035 : douta <= 12'h8A6 ;
		12'h036 : douta <= 12'h8A9 ;
		12'h037 : douta <= 12'h8AC ;
		12'h038 : douta <= 12'h8AF ;
		12'h039 : douta <= 12'h8B2 ;
		12'h03A : douta <= 12'h8B5 ;
		12'h03B : douta <= 12'h8B9 ;
		12'h03C : douta <= 12'h8BC ;
		12'h03D : douta <= 12'h8BF ;
		12'h03E : douta <= 12'h8C2 ;
		12'h03F : douta <= 12'h8C5 ;
		12'h040 : douta <= 12'h8C8 ;
		12'h041 : douta <= 12'h8CB ;
		12'h042 : douta <= 12'h8CE ;
		12'h043 : douta <= 12'h8D2 ;
		12'h044 : douta <= 12'h8D5 ;
		12'h045 : douta <= 12'h8D8 ;
		12'h046 : douta <= 12'h8DB ;
		12'h047 : douta <= 12'h8DE ;
		12'h048 : douta <= 12'h8E1 ;
		12'h049 : douta <= 12'h8E4 ;
		12'h04A : douta <= 12'h8E7 ;
		12'h04B : douta <= 12'h8EA ;
		12'h04C : douta <= 12'h8EE ;
		12'h04D : douta <= 12'h8F1 ;
		12'h04E : douta <= 12'h8F4 ;
		12'h04F : douta <= 12'h8F7 ;
		12'h050 : douta <= 12'h8FA ;
		12'h051 : douta <= 12'h8FD ;
		12'h052 : douta <= 12'h900 ;
		12'h053 : douta <= 12'h903 ;
		12'h054 : douta <= 12'h907 ;
		12'h055 : douta <= 12'h90A ;
		12'h056 : douta <= 12'h90D ;
		12'h057 : douta <= 12'h910 ;
		12'h058 : douta <= 12'h913 ;
		12'h059 : douta <= 12'h916 ;
		12'h05A : douta <= 12'h919 ;
		12'h05B : douta <= 12'h91C ;
		12'h05C : douta <= 12'h91F ;
		12'h05D : douta <= 12'h923 ;
		12'h05E : douta <= 12'h926 ;
		12'h05F : douta <= 12'h929 ;
		12'h060 : douta <= 12'h92C ;
		12'h061 : douta <= 12'h92F ;
		12'h062 : douta <= 12'h932 ;
		12'h063 : douta <= 12'h935 ;
		12'h064 : douta <= 12'h938 ;
		12'h065 : douta <= 12'h93B ;
		12'h066 : douta <= 12'h93E ;
		12'h067 : douta <= 12'h942 ;
		12'h068 : douta <= 12'h945 ;
		12'h069 : douta <= 12'h948 ;
		12'h06A : douta <= 12'h94B ;
		12'h06B : douta <= 12'h94E ;
		12'h06C : douta <= 12'h951 ;
		12'h06D : douta <= 12'h954 ;
		12'h06E : douta <= 12'h957 ;
		12'h06F : douta <= 12'h95A ;
		12'h070 : douta <= 12'h95D ;
		12'h071 : douta <= 12'h961 ;
		12'h072 : douta <= 12'h964 ;
		12'h073 : douta <= 12'h967 ;
		12'h074 : douta <= 12'h96A ;
		12'h075 : douta <= 12'h96D ;
		12'h076 : douta <= 12'h970 ;
		12'h077 : douta <= 12'h973 ;
		12'h078 : douta <= 12'h976 ;
		12'h079 : douta <= 12'h979 ;
		12'h07A : douta <= 12'h97C ;
		12'h07B : douta <= 12'h97F ;
		12'h07C : douta <= 12'h983 ;
		12'h07D : douta <= 12'h986 ;
		12'h07E : douta <= 12'h989 ;
		12'h07F : douta <= 12'h98C ;
		12'h080 : douta <= 12'h98F ;
		12'h081 : douta <= 12'h992 ;
		12'h082 : douta <= 12'h995 ;
		12'h083 : douta <= 12'h998 ;
		12'h084 : douta <= 12'h99B ;
		12'h085 : douta <= 12'h99E ;
		12'h086 : douta <= 12'h9A1 ;
		12'h087 : douta <= 12'h9A4 ;
		12'h088 : douta <= 12'h9A7 ;
		12'h089 : douta <= 12'h9AB ;
		12'h08A : douta <= 12'h9AE ;
		12'h08B : douta <= 12'h9B1 ;
		12'h08C : douta <= 12'h9B4 ;
		12'h08D : douta <= 12'h9B7 ;
		12'h08E : douta <= 12'h9BA ;
		12'h08F : douta <= 12'h9BD ;
		12'h090 : douta <= 12'h9C0 ;
		12'h091 : douta <= 12'h9C3 ;
		12'h092 : douta <= 12'h9C6 ;
		12'h093 : douta <= 12'h9C9 ;
		12'h094 : douta <= 12'h9CC ;
		12'h095 : douta <= 12'h9CF ;
		12'h096 : douta <= 12'h9D2 ;
		12'h097 : douta <= 12'h9D5 ;
		12'h098 : douta <= 12'h9D8 ;
		12'h099 : douta <= 12'h9DC ;
		12'h09A : douta <= 12'h9DF ;
		12'h09B : douta <= 12'h9E2 ;
		12'h09C : douta <= 12'h9E5 ;
		12'h09D : douta <= 12'h9E8 ;
		12'h09E : douta <= 12'h9EB ;
		12'h09F : douta <= 12'h9EE ;
		12'h0A0 : douta <= 12'h9F1 ;
		12'h0A1 : douta <= 12'h9F4 ;
		12'h0A2 : douta <= 12'h9F7 ;
		12'h0A3 : douta <= 12'h9FA ;
		12'h0A4 : douta <= 12'h9FD ;
		12'h0A5 : douta <= 12'hA00 ;
		12'h0A6 : douta <= 12'hA03 ;
		12'h0A7 : douta <= 12'hA06 ;
		12'h0A8 : douta <= 12'hA09 ;
		12'h0A9 : douta <= 12'hA0C ;
		12'h0AA : douta <= 12'hA0F ;
		12'h0AB : douta <= 12'hA12 ;
		12'h0AC : douta <= 12'hA15 ;
		12'h0AD : douta <= 12'hA18 ;
		12'h0AE : douta <= 12'hA1B ;
		12'h0AF : douta <= 12'hA1E ;
		12'h0B0 : douta <= 12'hA21 ;
		12'h0B1 : douta <= 12'hA24 ;
		12'h0B2 : douta <= 12'hA28 ;
		12'h0B3 : douta <= 12'hA2B ;
		12'h0B4 : douta <= 12'hA2E ;
		12'h0B5 : douta <= 12'hA31 ;
		12'h0B6 : douta <= 12'hA34 ;
		12'h0B7 : douta <= 12'hA37 ;
		12'h0B8 : douta <= 12'hA3A ;
		12'h0B9 : douta <= 12'hA3D ;
		12'h0BA : douta <= 12'hA40 ;
		12'h0BB : douta <= 12'hA43 ;
		12'h0BC : douta <= 12'hA46 ;
		12'h0BD : douta <= 12'hA49 ;
		12'h0BE : douta <= 12'hA4C ;
		12'h0BF : douta <= 12'hA4F ;
		12'h0C0 : douta <= 12'hA52 ;
		12'h0C1 : douta <= 12'hA55 ;
		12'h0C2 : douta <= 12'hA58 ;
		12'h0C3 : douta <= 12'hA5B ;
		12'h0C4 : douta <= 12'hA5E ;
		12'h0C5 : douta <= 12'hA61 ;
		12'h0C6 : douta <= 12'hA64 ;
		12'h0C7 : douta <= 12'hA67 ;
		12'h0C8 : douta <= 12'hA6A ;
		12'h0C9 : douta <= 12'hA6D ;
		12'h0CA : douta <= 12'hA70 ;
		12'h0CB : douta <= 12'hA73 ;
		12'h0CC : douta <= 12'hA76 ;
		12'h0CD : douta <= 12'hA79 ;
		12'h0CE : douta <= 12'hA7C ;
		12'h0CF : douta <= 12'hA7F ;
		12'h0D0 : douta <= 12'hA82 ;
		12'h0D1 : douta <= 12'hA85 ;
		12'h0D2 : douta <= 12'hA88 ;
		12'h0D3 : douta <= 12'hA8B ;
		12'h0D4 : douta <= 12'hA8E ;
		12'h0D5 : douta <= 12'hA90 ;
		12'h0D6 : douta <= 12'hA93 ;
		12'h0D7 : douta <= 12'hA96 ;
		12'h0D8 : douta <= 12'hA99 ;
		12'h0D9 : douta <= 12'hA9C ;
		12'h0DA : douta <= 12'hA9F ;
		12'h0DB : douta <= 12'hAA2 ;
		12'h0DC : douta <= 12'hAA5 ;
		12'h0DD : douta <= 12'hAA8 ;
		12'h0DE : douta <= 12'hAAB ;
		12'h0DF : douta <= 12'hAAE ;
		12'h0E0 : douta <= 12'hAB1 ;
		12'h0E1 : douta <= 12'hAB4 ;
		12'h0E2 : douta <= 12'hAB7 ;
		12'h0E3 : douta <= 12'hABA ;
		12'h0E4 : douta <= 12'hABD ;
		12'h0E5 : douta <= 12'hAC0 ;
		12'h0E6 : douta <= 12'hAC3 ;
		12'h0E7 : douta <= 12'hAC6 ;
		12'h0E8 : douta <= 12'hAC9 ;
		12'h0E9 : douta <= 12'hACC ;
		12'h0EA : douta <= 12'hACF ;
		12'h0EB : douta <= 12'hAD2 ;
		12'h0EC : douta <= 12'hAD4 ;
		12'h0ED : douta <= 12'hAD7 ;
		12'h0EE : douta <= 12'hADA ;
		12'h0EF : douta <= 12'hADD ;
		12'h0F0 : douta <= 12'hAE0 ;
		12'h0F1 : douta <= 12'hAE3 ;
		12'h0F2 : douta <= 12'hAE6 ;
		12'h0F3 : douta <= 12'hAE9 ;
		12'h0F4 : douta <= 12'hAEC ;
		12'h0F5 : douta <= 12'hAEF ;
		12'h0F6 : douta <= 12'hAF2 ;
		12'h0F7 : douta <= 12'hAF5 ;
		12'h0F8 : douta <= 12'hAF8 ;
		12'h0F9 : douta <= 12'hAFB ;
		12'h0FA : douta <= 12'hAFD ;
		12'h0FB : douta <= 12'hB00 ;
		12'h0FC : douta <= 12'hB03 ;
		12'h0FD : douta <= 12'hB06 ;
		12'h0FE : douta <= 12'hB09 ;
		12'h0FF : douta <= 12'hB0C ;
		12'h100 : douta <= 12'hB0F ;
		12'h101 : douta <= 12'hB12 ;
		12'h102 : douta <= 12'hB15 ;
		12'h103 : douta <= 12'hB18 ;
		12'h104 : douta <= 12'hB1A ;
		12'h105 : douta <= 12'hB1D ;
		12'h106 : douta <= 12'hB20 ;
		12'h107 : douta <= 12'hB23 ;
		12'h108 : douta <= 12'hB26 ;
		12'h109 : douta <= 12'hB29 ;
		12'h10A : douta <= 12'hB2C ;
		12'h10B : douta <= 12'hB2F ;
		12'h10C : douta <= 12'hB32 ;
		12'h10D : douta <= 12'hB34 ;
		12'h10E : douta <= 12'hB37 ;
		12'h10F : douta <= 12'hB3A ;
		12'h110 : douta <= 12'hB3D ;
		12'h111 : douta <= 12'hB40 ;
		12'h112 : douta <= 12'hB43 ;
		12'h113 : douta <= 12'hB46 ;
		12'h114 : douta <= 12'hB48 ;
		12'h115 : douta <= 12'hB4B ;
		12'h116 : douta <= 12'hB4E ;
		12'h117 : douta <= 12'hB51 ;
		12'h118 : douta <= 12'hB54 ;
		12'h119 : douta <= 12'hB57 ;
		12'h11A : douta <= 12'hB5A ;
		12'h11B : douta <= 12'hB5C ;
		12'h11C : douta <= 12'hB5F ;
		12'h11D : douta <= 12'hB62 ;
		12'h11E : douta <= 12'hB65 ;
		12'h11F : douta <= 12'hB68 ;
		12'h120 : douta <= 12'hB6B ;
		12'h121 : douta <= 12'hB6E ;
		12'h122 : douta <= 12'hB70 ;
		12'h123 : douta <= 12'hB73 ;
		12'h124 : douta <= 12'hB76 ;
		12'h125 : douta <= 12'hB79 ;
		12'h126 : douta <= 12'hB7C ;
		12'h127 : douta <= 12'hB7F ;
		12'h128 : douta <= 12'hB81 ;
		12'h129 : douta <= 12'hB84 ;
		12'h12A : douta <= 12'hB87 ;
		12'h12B : douta <= 12'hB8A ;
		12'h12C : douta <= 12'hB8D ;
		12'h12D : douta <= 12'hB8F ;
		12'h12E : douta <= 12'hB92 ;
		12'h12F : douta <= 12'hB95 ;
		12'h130 : douta <= 12'hB98 ;
		12'h131 : douta <= 12'hB9B ;
		12'h132 : douta <= 12'hB9D ;
		12'h133 : douta <= 12'hBA0 ;
		12'h134 : douta <= 12'hBA3 ;
		12'h135 : douta <= 12'hBA6 ;
		12'h136 : douta <= 12'hBA9 ;
		12'h137 : douta <= 12'hBAB ;
		12'h138 : douta <= 12'hBAE ;
		12'h139 : douta <= 12'hBB1 ;
		12'h13A : douta <= 12'hBB4 ;
		12'h13B : douta <= 12'hBB7 ;
		12'h13C : douta <= 12'hBB9 ;
		12'h13D : douta <= 12'hBBC ;
		12'h13E : douta <= 12'hBBF ;
		12'h13F : douta <= 12'hBC2 ;
		12'h140 : douta <= 12'hBC4 ;
		12'h141 : douta <= 12'hBC7 ;
		12'h142 : douta <= 12'hBCA ;
		12'h143 : douta <= 12'hBCD ;
		12'h144 : douta <= 12'hBD0 ;
		12'h145 : douta <= 12'hBD2 ;
		12'h146 : douta <= 12'hBD5 ;
		12'h147 : douta <= 12'hBD8 ;
		12'h148 : douta <= 12'hBDB ;
		12'h149 : douta <= 12'hBDD ;
		12'h14A : douta <= 12'hBE0 ;
		12'h14B : douta <= 12'hBE3 ;
		12'h14C : douta <= 12'hBE6 ;
		12'h14D : douta <= 12'hBE8 ;
		12'h14E : douta <= 12'hBEB ;
		12'h14F : douta <= 12'hBEE ;
		12'h150 : douta <= 12'hBF0 ;
		12'h151 : douta <= 12'hBF3 ;
		12'h152 : douta <= 12'hBF6 ;
		12'h153 : douta <= 12'hBF9 ;
		12'h154 : douta <= 12'hBFB ;
		12'h155 : douta <= 12'hBFE ;
		12'h156 : douta <= 12'hC01 ;
		12'h157 : douta <= 12'hC04 ;
		12'h158 : douta <= 12'hC06 ;
		12'h159 : douta <= 12'hC09 ;
		12'h15A : douta <= 12'hC0C ;
		12'h15B : douta <= 12'hC0E ;
		12'h15C : douta <= 12'hC11 ;
		12'h15D : douta <= 12'hC14 ;
		12'h15E : douta <= 12'hC16 ;
		12'h15F : douta <= 12'hC19 ;
		12'h160 : douta <= 12'hC1C ;
		12'h161 : douta <= 12'hC1F ;
		12'h162 : douta <= 12'hC21 ;
		12'h163 : douta <= 12'hC24 ;
		12'h164 : douta <= 12'hC27 ;
		12'h165 : douta <= 12'hC29 ;
		12'h166 : douta <= 12'hC2C ;
		12'h167 : douta <= 12'hC2F ;
		12'h168 : douta <= 12'hC31 ;
		12'h169 : douta <= 12'hC34 ;
		12'h16A : douta <= 12'hC37 ;
		12'h16B : douta <= 12'hC39 ;
		12'h16C : douta <= 12'hC3C ;
		12'h16D : douta <= 12'hC3F ;
		12'h16E : douta <= 12'hC41 ;
		12'h16F : douta <= 12'hC44 ;
		12'h170 : douta <= 12'hC47 ;
		12'h171 : douta <= 12'hC49 ;
		12'h172 : douta <= 12'hC4C ;
		12'h173 : douta <= 12'hC4F ;
		12'h174 : douta <= 12'hC51 ;
		12'h175 : douta <= 12'hC54 ;
		12'h176 : douta <= 12'hC57 ;
		12'h177 : douta <= 12'hC59 ;
		12'h178 : douta <= 12'hC5C ;
		12'h179 : douta <= 12'hC5E ;
		12'h17A : douta <= 12'hC61 ;
		12'h17B : douta <= 12'hC64 ;
		12'h17C : douta <= 12'hC66 ;
		12'h17D : douta <= 12'hC69 ;
		12'h17E : douta <= 12'hC6C ;
		12'h17F : douta <= 12'hC6E ;
		12'h180 : douta <= 12'hC71 ;
		12'h181 : douta <= 12'hC73 ;
		12'h182 : douta <= 12'hC76 ;
		12'h183 : douta <= 12'hC79 ;
		12'h184 : douta <= 12'hC7B ;
		12'h185 : douta <= 12'hC7E ;
		12'h186 : douta <= 12'hC80 ;
		12'h187 : douta <= 12'hC83 ;
		12'h188 : douta <= 12'hC86 ;
		12'h189 : douta <= 12'hC88 ;
		12'h18A : douta <= 12'hC8B ;
		12'h18B : douta <= 12'hC8D ;
		12'h18C : douta <= 12'hC90 ;
		12'h18D : douta <= 12'hC92 ;
		12'h18E : douta <= 12'hC95 ;
		12'h18F : douta <= 12'hC98 ;
		12'h190 : douta <= 12'hC9A ;
		12'h191 : douta <= 12'hC9D ;
		12'h192 : douta <= 12'hC9F ;
		12'h193 : douta <= 12'hCA2 ;
		12'h194 : douta <= 12'hCA4 ;
		12'h195 : douta <= 12'hCA7 ;
		12'h196 : douta <= 12'hCAA ;
		12'h197 : douta <= 12'hCAC ;
		12'h198 : douta <= 12'hCAF ;
		12'h199 : douta <= 12'hCB1 ;
		12'h19A : douta <= 12'hCB4 ;
		12'h19B : douta <= 12'hCB6 ;
		12'h19C : douta <= 12'hCB9 ;
		12'h19D : douta <= 12'hCBB ;
		12'h19E : douta <= 12'hCBE ;
		12'h19F : douta <= 12'hCC0 ;
		12'h1A0 : douta <= 12'hCC3 ;
		12'h1A1 : douta <= 12'hCC5 ;
		12'h1A2 : douta <= 12'hCC8 ;
		12'h1A3 : douta <= 12'hCCA ;
		12'h1A4 : douta <= 12'hCCD ;
		12'h1A5 : douta <= 12'hCCF ;
		12'h1A6 : douta <= 12'hCD2 ;
		12'h1A7 : douta <= 12'hCD4 ;
		12'h1A8 : douta <= 12'hCD7 ;
		12'h1A9 : douta <= 12'hCD9 ;
		12'h1AA : douta <= 12'hCDC ;
		12'h1AB : douta <= 12'hCDE ;
		12'h1AC : douta <= 12'hCE1 ;
		12'h1AD : douta <= 12'hCE3 ;
		12'h1AE : douta <= 12'hCE6 ;
		12'h1AF : douta <= 12'hCE8 ;
		12'h1B0 : douta <= 12'hCEB ;
		12'h1B1 : douta <= 12'hCED ;
		12'h1B2 : douta <= 12'hCF0 ;
		12'h1B3 : douta <= 12'hCF2 ;
		12'h1B4 : douta <= 12'hCF5 ;
		12'h1B5 : douta <= 12'hCF7 ;
		12'h1B6 : douta <= 12'hCFA ;
		12'h1B7 : douta <= 12'hCFC ;
		12'h1B8 : douta <= 12'hCFF ;
		12'h1B9 : douta <= 12'hD01 ;
		12'h1BA : douta <= 12'hD03 ;
		12'h1BB : douta <= 12'hD06 ;
		12'h1BC : douta <= 12'hD08 ;
		12'h1BD : douta <= 12'hD0B ;
		12'h1BE : douta <= 12'hD0D ;
		12'h1BF : douta <= 12'hD10 ;
		12'h1C0 : douta <= 12'hD12 ;
		12'h1C1 : douta <= 12'hD15 ;
		12'h1C2 : douta <= 12'hD17 ;
		12'h1C3 : douta <= 12'hD19 ;
		12'h1C4 : douta <= 12'hD1C ;
		12'h1C5 : douta <= 12'hD1E ;
		12'h1C6 : douta <= 12'hD21 ;
		12'h1C7 : douta <= 12'hD23 ;
		12'h1C8 : douta <= 12'hD25 ;
		12'h1C9 : douta <= 12'hD28 ;
		12'h1CA : douta <= 12'hD2A ;
		12'h1CB : douta <= 12'hD2D ;
		12'h1CC : douta <= 12'hD2F ;
		12'h1CD : douta <= 12'hD31 ;
		12'h1CE : douta <= 12'hD34 ;
		12'h1CF : douta <= 12'hD36 ;
		12'h1D0 : douta <= 12'hD39 ;
		12'h1D1 : douta <= 12'hD3B ;
		12'h1D2 : douta <= 12'hD3D ;
		12'h1D3 : douta <= 12'hD40 ;
		12'h1D4 : douta <= 12'hD42 ;
		12'h1D5 : douta <= 12'hD44 ;
		12'h1D6 : douta <= 12'hD47 ;
		12'h1D7 : douta <= 12'hD49 ;
		12'h1D8 : douta <= 12'hD4B ;
		12'h1D9 : douta <= 12'hD4E ;
		12'h1DA : douta <= 12'hD50 ;
		12'h1DB : douta <= 12'hD53 ;
		12'h1DC : douta <= 12'hD55 ;
		12'h1DD : douta <= 12'hD57 ;
		12'h1DE : douta <= 12'hD5A ;
		12'h1DF : douta <= 12'hD5C ;
		12'h1E0 : douta <= 12'hD5E ;
		12'h1E1 : douta <= 12'hD61 ;
		12'h1E2 : douta <= 12'hD63 ;
		12'h1E3 : douta <= 12'hD65 ;
		12'h1E4 : douta <= 12'hD67 ;
		12'h1E5 : douta <= 12'hD6A ;
		12'h1E6 : douta <= 12'hD6C ;
		12'h1E7 : douta <= 12'hD6E ;
		12'h1E8 : douta <= 12'hD71 ;
		12'h1E9 : douta <= 12'hD73 ;
		12'h1EA : douta <= 12'hD75 ;
		12'h1EB : douta <= 12'hD78 ;
		12'h1EC : douta <= 12'hD7A ;
		12'h1ED : douta <= 12'hD7C ;
		12'h1EE : douta <= 12'hD7E ;
		12'h1EF : douta <= 12'hD81 ;
		12'h1F0 : douta <= 12'hD83 ;
		12'h1F1 : douta <= 12'hD85 ;
		12'h1F2 : douta <= 12'hD88 ;
		12'h1F3 : douta <= 12'hD8A ;
		12'h1F4 : douta <= 12'hD8C ;
		12'h1F5 : douta <= 12'hD8E ;
		12'h1F6 : douta <= 12'hD91 ;
		12'h1F7 : douta <= 12'hD93 ;
		12'h1F8 : douta <= 12'hD95 ;
		12'h1F9 : douta <= 12'hD97 ;
		12'h1FA : douta <= 12'hD9A ;
		12'h1FB : douta <= 12'hD9C ;
		12'h1FC : douta <= 12'hD9E ;
		12'h1FD : douta <= 12'hDA0 ;
		12'h1FE : douta <= 12'hDA3 ;
		12'h1FF : douta <= 12'hDA5 ;
		12'h200 : douta <= 12'hDA7 ;
		12'h201 : douta <= 12'hDA9 ;
		12'h202 : douta <= 12'hDAB ;
		12'h203 : douta <= 12'hDAE ;
		12'h204 : douta <= 12'hDB0 ;
		12'h205 : douta <= 12'hDB2 ;
		12'h206 : douta <= 12'hDB4 ;
		12'h207 : douta <= 12'hDB6 ;
		12'h208 : douta <= 12'hDB9 ;
		12'h209 : douta <= 12'hDBB ;
		12'h20A : douta <= 12'hDBD ;
		12'h20B : douta <= 12'hDBF ;
		12'h20C : douta <= 12'hDC1 ;
		12'h20D : douta <= 12'hDC4 ;
		12'h20E : douta <= 12'hDC6 ;
		12'h20F : douta <= 12'hDC8 ;
		12'h210 : douta <= 12'hDCA ;
		12'h211 : douta <= 12'hDCC ;
		12'h212 : douta <= 12'hDCE ;
		12'h213 : douta <= 12'hDD1 ;
		12'h214 : douta <= 12'hDD3 ;
		12'h215 : douta <= 12'hDD5 ;
		12'h216 : douta <= 12'hDD7 ;
		12'h217 : douta <= 12'hDD9 ;
		12'h218 : douta <= 12'hDDB ;
		12'h219 : douta <= 12'hDDD ;
		12'h21A : douta <= 12'hDE0 ;
		12'h21B : douta <= 12'hDE2 ;
		12'h21C : douta <= 12'hDE4 ;
		12'h21D : douta <= 12'hDE6 ;
		12'h21E : douta <= 12'hDE8 ;
		12'h21F : douta <= 12'hDEA ;
		12'h220 : douta <= 12'hDEC ;
		12'h221 : douta <= 12'hDEE ;
		12'h222 : douta <= 12'hDF0 ;
		12'h223 : douta <= 12'hDF3 ;
		12'h224 : douta <= 12'hDF5 ;
		12'h225 : douta <= 12'hDF7 ;
		12'h226 : douta <= 12'hDF9 ;
		12'h227 : douta <= 12'hDFB ;
		12'h228 : douta <= 12'hDFD ;
		12'h229 : douta <= 12'hDFF ;
		12'h22A : douta <= 12'hE01 ;
		12'h22B : douta <= 12'hE03 ;
		12'h22C : douta <= 12'hE05 ;
		12'h22D : douta <= 12'hE07 ;
		12'h22E : douta <= 12'hE09 ;
		12'h22F : douta <= 12'hE0B ;
		12'h230 : douta <= 12'hE0E ;
		12'h231 : douta <= 12'hE10 ;
		12'h232 : douta <= 12'hE12 ;
		12'h233 : douta <= 12'hE14 ;
		12'h234 : douta <= 12'hE16 ;
		12'h235 : douta <= 12'hE18 ;
		12'h236 : douta <= 12'hE1A ;
		12'h237 : douta <= 12'hE1C ;
		12'h238 : douta <= 12'hE1E ;
		12'h239 : douta <= 12'hE20 ;
		12'h23A : douta <= 12'hE22 ;
		12'h23B : douta <= 12'hE24 ;
		12'h23C : douta <= 12'hE26 ;
		12'h23D : douta <= 12'hE28 ;
		12'h23E : douta <= 12'hE2A ;
		12'h23F : douta <= 12'hE2C ;
		12'h240 : douta <= 12'hE2E ;
		12'h241 : douta <= 12'hE30 ;
		12'h242 : douta <= 12'hE32 ;
		12'h243 : douta <= 12'hE34 ;
		12'h244 : douta <= 12'hE36 ;
		12'h245 : douta <= 12'hE38 ;
		12'h246 : douta <= 12'hE3A ;
		12'h247 : douta <= 12'hE3C ;
		12'h248 : douta <= 12'hE3E ;
		12'h249 : douta <= 12'hE40 ;
		12'h24A : douta <= 12'hE42 ;
		12'h24B : douta <= 12'hE44 ;
		12'h24C : douta <= 12'hE45 ;
		12'h24D : douta <= 12'hE47 ;
		12'h24E : douta <= 12'hE49 ;
		12'h24F : douta <= 12'hE4B ;
		12'h250 : douta <= 12'hE4D ;
		12'h251 : douta <= 12'hE4F ;
		12'h252 : douta <= 12'hE51 ;
		12'h253 : douta <= 12'hE53 ;
		12'h254 : douta <= 12'hE55 ;
		12'h255 : douta <= 12'hE57 ;
		12'h256 : douta <= 12'hE59 ;
		12'h257 : douta <= 12'hE5B ;
		12'h258 : douta <= 12'hE5D ;
		12'h259 : douta <= 12'hE5E ;
		12'h25A : douta <= 12'hE60 ;
		12'h25B : douta <= 12'hE62 ;
		12'h25C : douta <= 12'hE64 ;
		12'h25D : douta <= 12'hE66 ;
		12'h25E : douta <= 12'hE68 ;
		12'h25F : douta <= 12'hE6A ;
		12'h260 : douta <= 12'hE6C ;
		12'h261 : douta <= 12'hE6E ;
		12'h262 : douta <= 12'hE6F ;
		12'h263 : douta <= 12'hE71 ;
		12'h264 : douta <= 12'hE73 ;
		12'h265 : douta <= 12'hE75 ;
		12'h266 : douta <= 12'hE77 ;
		12'h267 : douta <= 12'hE79 ;
		12'h268 : douta <= 12'hE7B ;
		12'h269 : douta <= 12'hE7C ;
		12'h26A : douta <= 12'hE7E ;
		12'h26B : douta <= 12'hE80 ;
		12'h26C : douta <= 12'hE82 ;
		12'h26D : douta <= 12'hE84 ;
		12'h26E : douta <= 12'hE85 ;
		12'h26F : douta <= 12'hE87 ;
		12'h270 : douta <= 12'hE89 ;
		12'h271 : douta <= 12'hE8B ;
		12'h272 : douta <= 12'hE8D ;
		12'h273 : douta <= 12'hE8F ;
		12'h274 : douta <= 12'hE90 ;
		12'h275 : douta <= 12'hE92 ;
		12'h276 : douta <= 12'hE94 ;
		12'h277 : douta <= 12'hE96 ;
		12'h278 : douta <= 12'hE97 ;
		12'h279 : douta <= 12'hE99 ;
		12'h27A : douta <= 12'hE9B ;
		12'h27B : douta <= 12'hE9D ;
		12'h27C : douta <= 12'hE9F ;
		12'h27D : douta <= 12'hEA0 ;
		12'h27E : douta <= 12'hEA2 ;
		12'h27F : douta <= 12'hEA4 ;
		12'h280 : douta <= 12'hEA6 ;
		12'h281 : douta <= 12'hEA7 ;
		12'h282 : douta <= 12'hEA9 ;
		12'h283 : douta <= 12'hEAB ;
		12'h284 : douta <= 12'hEAC ;
		12'h285 : douta <= 12'hEAE ;
		12'h286 : douta <= 12'hEB0 ;
		12'h287 : douta <= 12'hEB2 ;
		12'h288 : douta <= 12'hEB3 ;
		12'h289 : douta <= 12'hEB5 ;
		12'h28A : douta <= 12'hEB7 ;
		12'h28B : douta <= 12'hEB8 ;
		12'h28C : douta <= 12'hEBA ;
		12'h28D : douta <= 12'hEBC ;
		12'h28E : douta <= 12'hEBE ;
		12'h28F : douta <= 12'hEBF ;
		12'h290 : douta <= 12'hEC1 ;
		12'h291 : douta <= 12'hEC3 ;
		12'h292 : douta <= 12'hEC4 ;
		12'h293 : douta <= 12'hEC6 ;
		12'h294 : douta <= 12'hEC8 ;
		12'h295 : douta <= 12'hEC9 ;
		12'h296 : douta <= 12'hECB ;
		12'h297 : douta <= 12'hECD ;
		12'h298 : douta <= 12'hECE ;
		12'h299 : douta <= 12'hED0 ;
		12'h29A : douta <= 12'hED2 ;
		12'h29B : douta <= 12'hED3 ;
		12'h29C : douta <= 12'hED5 ;
		12'h29D : douta <= 12'hED6 ;
		12'h29E : douta <= 12'hED8 ;
		12'h29F : douta <= 12'hEDA ;
		12'h2A0 : douta <= 12'hEDB ;
		12'h2A1 : douta <= 12'hEDD ;
		12'h2A2 : douta <= 12'hEDE ;
		12'h2A3 : douta <= 12'hEE0 ;
		12'h2A4 : douta <= 12'hEE2 ;
		12'h2A5 : douta <= 12'hEE3 ;
		12'h2A6 : douta <= 12'hEE5 ;
		12'h2A7 : douta <= 12'hEE6 ;
		12'h2A8 : douta <= 12'hEE8 ;
		12'h2A9 : douta <= 12'hEEA ;
		12'h2AA : douta <= 12'hEEB ;
		12'h2AB : douta <= 12'hEED ;
		12'h2AC : douta <= 12'hEEE ;
		12'h2AD : douta <= 12'hEF0 ;
		12'h2AE : douta <= 12'hEF1 ;
		12'h2AF : douta <= 12'hEF3 ;
		12'h2B0 : douta <= 12'hEF5 ;
		12'h2B1 : douta <= 12'hEF6 ;
		12'h2B2 : douta <= 12'hEF8 ;
		12'h2B3 : douta <= 12'hEF9 ;
		12'h2B4 : douta <= 12'hEFB ;
		12'h2B5 : douta <= 12'hEFC ;
		12'h2B6 : douta <= 12'hEFE ;
		12'h2B7 : douta <= 12'hEFF ;
		12'h2B8 : douta <= 12'hF01 ;
		12'h2B9 : douta <= 12'hF02 ;
		12'h2BA : douta <= 12'hF04 ;
		12'h2BB : douta <= 12'hF05 ;
		12'h2BC : douta <= 12'hF07 ;
		12'h2BD : douta <= 12'hF08 ;
		12'h2BE : douta <= 12'hF0A ;
		12'h2BF : douta <= 12'hF0B ;
		12'h2C0 : douta <= 12'hF0D ;
		12'h2C1 : douta <= 12'hF0E ;
		12'h2C2 : douta <= 12'hF10 ;
		12'h2C3 : douta <= 12'hF11 ;
		12'h2C4 : douta <= 12'hF13 ;
		12'h2C5 : douta <= 12'hF14 ;
		12'h2C6 : douta <= 12'hF16 ;
		12'h2C7 : douta <= 12'hF17 ;
		12'h2C8 : douta <= 12'hF18 ;
		12'h2C9 : douta <= 12'hF1A ;
		12'h2CA : douta <= 12'hF1B ;
		12'h2CB : douta <= 12'hF1D ;
		12'h2CC : douta <= 12'hF1E ;
		12'h2CD : douta <= 12'hF20 ;
		12'h2CE : douta <= 12'hF21 ;
		12'h2CF : douta <= 12'hF23 ;
		12'h2D0 : douta <= 12'hF24 ;
		12'h2D1 : douta <= 12'hF25 ;
		12'h2D2 : douta <= 12'hF27 ;
		12'h2D3 : douta <= 12'hF28 ;
		12'h2D4 : douta <= 12'hF2A ;
		12'h2D5 : douta <= 12'hF2B ;
		12'h2D6 : douta <= 12'hF2C ;
		12'h2D7 : douta <= 12'hF2E ;
		12'h2D8 : douta <= 12'hF2F ;
		12'h2D9 : douta <= 12'hF30 ;
		12'h2DA : douta <= 12'hF32 ;
		12'h2DB : douta <= 12'hF33 ;
		12'h2DC : douta <= 12'hF35 ;
		12'h2DD : douta <= 12'hF36 ;
		12'h2DE : douta <= 12'hF37 ;
		12'h2DF : douta <= 12'hF39 ;
		12'h2E0 : douta <= 12'hF3A ;
		12'h2E1 : douta <= 12'hF3B ;
		12'h2E2 : douta <= 12'hF3D ;
		12'h2E3 : douta <= 12'hF3E ;
		12'h2E4 : douta <= 12'hF3F ;
		12'h2E5 : douta <= 12'hF41 ;
		12'h2E6 : douta <= 12'hF42 ;
		12'h2E7 : douta <= 12'hF43 ;
		12'h2E8 : douta <= 12'hF45 ;
		12'h2E9 : douta <= 12'hF46 ;
		12'h2EA : douta <= 12'hF47 ;
		12'h2EB : douta <= 12'hF48 ;
		12'h2EC : douta <= 12'hF4A ;
		12'h2ED : douta <= 12'hF4B ;
		12'h2EE : douta <= 12'hF4C ;
		12'h2EF : douta <= 12'hF4E ;
		12'h2F0 : douta <= 12'hF4F ;
		12'h2F1 : douta <= 12'hF50 ;
		12'h2F2 : douta <= 12'hF51 ;
		12'h2F3 : douta <= 12'hF53 ;
		12'h2F4 : douta <= 12'hF54 ;
		12'h2F5 : douta <= 12'hF55 ;
		12'h2F6 : douta <= 12'hF56 ;
		12'h2F7 : douta <= 12'hF58 ;
		12'h2F8 : douta <= 12'hF59 ;
		12'h2F9 : douta <= 12'hF5A ;
		12'h2FA : douta <= 12'hF5B ;
		12'h2FB : douta <= 12'hF5D ;
		12'h2FC : douta <= 12'hF5E ;
		12'h2FD : douta <= 12'hF5F ;
		12'h2FE : douta <= 12'hF60 ;
		12'h2FF : douta <= 12'hF61 ;
		12'h300 : douta <= 12'hF63 ;
		12'h301 : douta <= 12'hF64 ;
		12'h302 : douta <= 12'hF65 ;
		12'h303 : douta <= 12'hF66 ;
		12'h304 : douta <= 12'hF67 ;
		12'h305 : douta <= 12'hF69 ;
		12'h306 : douta <= 12'hF6A ;
		12'h307 : douta <= 12'hF6B ;
		12'h308 : douta <= 12'hF6C ;
		12'h309 : douta <= 12'hF6D ;
		12'h30A : douta <= 12'hF6E ;
		12'h30B : douta <= 12'hF70 ;
		12'h30C : douta <= 12'hF71 ;
		12'h30D : douta <= 12'hF72 ;
		12'h30E : douta <= 12'hF73 ;
		12'h30F : douta <= 12'hF74 ;
		12'h310 : douta <= 12'hF75 ;
		12'h311 : douta <= 12'hF76 ;
		12'h312 : douta <= 12'hF78 ;
		12'h313 : douta <= 12'hF79 ;
		12'h314 : douta <= 12'hF7A ;
		12'h315 : douta <= 12'hF7B ;
		12'h316 : douta <= 12'hF7C ;
		12'h317 : douta <= 12'hF7D ;
		12'h318 : douta <= 12'hF7E ;
		12'h319 : douta <= 12'hF7F ;
		12'h31A : douta <= 12'hF80 ;
		12'h31B : douta <= 12'hF81 ;
		12'h31C : douta <= 12'hF83 ;
		12'h31D : douta <= 12'hF84 ;
		12'h31E : douta <= 12'hF85 ;
		12'h31F : douta <= 12'hF86 ;
		12'h320 : douta <= 12'hF87 ;
		12'h321 : douta <= 12'hF88 ;
		12'h322 : douta <= 12'hF89 ;
		12'h323 : douta <= 12'hF8A ;
		12'h324 : douta <= 12'hF8B ;
		12'h325 : douta <= 12'hF8C ;
		12'h326 : douta <= 12'hF8D ;
		12'h327 : douta <= 12'hF8E ;
		12'h328 : douta <= 12'hF8F ;
		12'h329 : douta <= 12'hF90 ;
		12'h32A : douta <= 12'hF91 ;
		12'h32B : douta <= 12'hF92 ;
		12'h32C : douta <= 12'hF93 ;
		12'h32D : douta <= 12'hF94 ;
		12'h32E : douta <= 12'hF95 ;
		12'h32F : douta <= 12'hF96 ;
		12'h330 : douta <= 12'hF97 ;
		12'h331 : douta <= 12'hF98 ;
		12'h332 : douta <= 12'hF99 ;
		12'h333 : douta <= 12'hF9A ;
		12'h334 : douta <= 12'hF9B ;
		12'h335 : douta <= 12'hF9C ;
		12'h336 : douta <= 12'hF9D ;
		12'h337 : douta <= 12'hF9E ;
		12'h338 : douta <= 12'hF9F ;
		12'h339 : douta <= 12'hFA0 ;
		12'h33A : douta <= 12'hFA1 ;
		12'h33B : douta <= 12'hFA2 ;
		12'h33C : douta <= 12'hFA3 ;
		12'h33D : douta <= 12'hFA4 ;
		12'h33E : douta <= 12'hFA5 ;
		12'h33F : douta <= 12'hFA5 ;
		12'h340 : douta <= 12'hFA6 ;
		12'h341 : douta <= 12'hFA7 ;
		12'h342 : douta <= 12'hFA8 ;
		12'h343 : douta <= 12'hFA9 ;
		12'h344 : douta <= 12'hFAA ;
		12'h345 : douta <= 12'hFAB ;
		12'h346 : douta <= 12'hFAC ;
		12'h347 : douta <= 12'hFAD ;
		12'h348 : douta <= 12'hFAE ;
		12'h349 : douta <= 12'hFAE ;
		12'h34A : douta <= 12'hFAF ;
		12'h34B : douta <= 12'hFB0 ;
		12'h34C : douta <= 12'hFB1 ;
		12'h34D : douta <= 12'hFB2 ;
		12'h34E : douta <= 12'hFB3 ;
		12'h34F : douta <= 12'hFB4 ;
		12'h350 : douta <= 12'hFB4 ;
		12'h351 : douta <= 12'hFB5 ;
		12'h352 : douta <= 12'hFB6 ;
		12'h353 : douta <= 12'hFB7 ;
		12'h354 : douta <= 12'hFB8 ;
		12'h355 : douta <= 12'hFB8 ;
		12'h356 : douta <= 12'hFB9 ;
		12'h357 : douta <= 12'hFBA ;
		12'h358 : douta <= 12'hFBB ;
		12'h359 : douta <= 12'hFBC ;
		12'h35A : douta <= 12'hFBC ;
		12'h35B : douta <= 12'hFBD ;
		12'h35C : douta <= 12'hFBE ;
		12'h35D : douta <= 12'hFBF ;
		12'h35E : douta <= 12'hFC0 ;
		12'h35F : douta <= 12'hFC0 ;
		12'h360 : douta <= 12'hFC1 ;
		12'h361 : douta <= 12'hFC2 ;
		12'h362 : douta <= 12'hFC3 ;
		12'h363 : douta <= 12'hFC3 ;
		12'h364 : douta <= 12'hFC4 ;
		12'h365 : douta <= 12'hFC5 ;
		12'h366 : douta <= 12'hFC6 ;
		12'h367 : douta <= 12'hFC6 ;
		12'h368 : douta <= 12'hFC7 ;
		12'h369 : douta <= 12'hFC8 ;
		12'h36A : douta <= 12'hFC9 ;
		12'h36B : douta <= 12'hFC9 ;
		12'h36C : douta <= 12'hFCA ;
		12'h36D : douta <= 12'hFCB ;
		12'h36E : douta <= 12'hFCB ;
		12'h36F : douta <= 12'hFCC ;
		12'h370 : douta <= 12'hFCD ;
		12'h371 : douta <= 12'hFCD ;
		12'h372 : douta <= 12'hFCE ;
		12'h373 : douta <= 12'hFCF ;
		12'h374 : douta <= 12'hFCF ;
		12'h375 : douta <= 12'hFD0 ;
		12'h376 : douta <= 12'hFD1 ;
		12'h377 : douta <= 12'hFD1 ;
		12'h378 : douta <= 12'hFD2 ;
		12'h379 : douta <= 12'hFD3 ;
		12'h37A : douta <= 12'hFD3 ;
		12'h37B : douta <= 12'hFD4 ;
		12'h37C : douta <= 12'hFD5 ;
		12'h37D : douta <= 12'hFD5 ;
		12'h37E : douta <= 12'hFD6 ;
		12'h37F : douta <= 12'hFD7 ;
		12'h380 : douta <= 12'hFD7 ;
		12'h381 : douta <= 12'hFD8 ;
		12'h382 : douta <= 12'hFD8 ;
		12'h383 : douta <= 12'hFD9 ;
		12'h384 : douta <= 12'hFDA ;
		12'h385 : douta <= 12'hFDA ;
		12'h386 : douta <= 12'hFDB ;
		12'h387 : douta <= 12'hFDB ;
		12'h388 : douta <= 12'hFDC ;
		12'h389 : douta <= 12'hFDC ;
		12'h38A : douta <= 12'hFDD ;
		12'h38B : douta <= 12'hFDE ;
		12'h38C : douta <= 12'hFDE ;
		12'h38D : douta <= 12'hFDF ;
		12'h38E : douta <= 12'hFDF ;
		12'h38F : douta <= 12'hFE0 ;
		12'h390 : douta <= 12'hFE0 ;
		12'h391 : douta <= 12'hFE1 ;
		12'h392 : douta <= 12'hFE1 ;
		12'h393 : douta <= 12'hFE2 ;
		12'h394 : douta <= 12'hFE2 ;
		12'h395 : douta <= 12'hFE3 ;
		12'h396 : douta <= 12'hFE3 ;
		12'h397 : douta <= 12'hFE4 ;
		12'h398 : douta <= 12'hFE5 ;
		12'h399 : douta <= 12'hFE5 ;
		12'h39A : douta <= 12'hFE5 ;
		12'h39B : douta <= 12'hFE6 ;
		12'h39C : douta <= 12'hFE6 ;
		12'h39D : douta <= 12'hFE7 ;
		12'h39E : douta <= 12'hFE7 ;
		12'h39F : douta <= 12'hFE8 ;
		12'h3A0 : douta <= 12'hFE8 ;
		12'h3A1 : douta <= 12'hFE9 ;
		12'h3A2 : douta <= 12'hFE9 ;
		12'h3A3 : douta <= 12'hFEA ;
		12'h3A4 : douta <= 12'hFEA ;
		12'h3A5 : douta <= 12'hFEB ;
		12'h3A6 : douta <= 12'hFEB ;
		12'h3A7 : douta <= 12'hFEB ;
		12'h3A8 : douta <= 12'hFEC ;
		12'h3A9 : douta <= 12'hFEC ;
		12'h3AA : douta <= 12'hFED ;
		12'h3AB : douta <= 12'hFED ;
		12'h3AC : douta <= 12'hFEE ;
		12'h3AD : douta <= 12'hFEE ;
		12'h3AE : douta <= 12'hFEE ;
		12'h3AF : douta <= 12'hFEF ;
		12'h3B0 : douta <= 12'hFEF ;
		12'h3B1 : douta <= 12'hFEF ;
		12'h3B2 : douta <= 12'hFF0 ;
		12'h3B3 : douta <= 12'hFF0 ;
		12'h3B4 : douta <= 12'hFF1 ;
		12'h3B5 : douta <= 12'hFF1 ;
		12'h3B6 : douta <= 12'hFF1 ;
		12'h3B7 : douta <= 12'hFF2 ;
		12'h3B8 : douta <= 12'hFF2 ;
		12'h3B9 : douta <= 12'hFF2 ;
		12'h3BA : douta <= 12'hFF3 ;
		12'h3BB : douta <= 12'hFF3 ;
		12'h3BC : douta <= 12'hFF3 ;
		12'h3BD : douta <= 12'hFF4 ;
		12'h3BE : douta <= 12'hFF4 ;
		12'h3BF : douta <= 12'hFF4 ;
		12'h3C0 : douta <= 12'hFF5 ;
		12'h3C1 : douta <= 12'hFF5 ;
		12'h3C2 : douta <= 12'hFF5 ;
		12'h3C3 : douta <= 12'hFF6 ;
		12'h3C4 : douta <= 12'hFF6 ;
		12'h3C5 : douta <= 12'hFF6 ;
		12'h3C6 : douta <= 12'hFF6 ;
		12'h3C7 : douta <= 12'hFF7 ;
		12'h3C8 : douta <= 12'hFF7 ;
		12'h3C9 : douta <= 12'hFF7 ;
		12'h3CA : douta <= 12'hFF7 ;
		12'h3CB : douta <= 12'hFF8 ;
		12'h3CC : douta <= 12'hFF8 ;
		12'h3CD : douta <= 12'hFF8 ;
		12'h3CE : douta <= 12'hFF8 ;
		12'h3CF : douta <= 12'hFF9 ;
		12'h3D0 : douta <= 12'hFF9 ;
		12'h3D1 : douta <= 12'hFF9 ;
		12'h3D2 : douta <= 12'hFF9 ;
		12'h3D3 : douta <= 12'hFFA ;
		12'h3D4 : douta <= 12'hFFA ;
		12'h3D5 : douta <= 12'hFFA ;
		12'h3D6 : douta <= 12'hFFA ;
		12'h3D7 : douta <= 12'hFFA ;
		12'h3D8 : douta <= 12'hFFB ;
		12'h3D9 : douta <= 12'hFFB ;
		12'h3DA : douta <= 12'hFFB ;
		12'h3DB : douta <= 12'hFFB ;
		12'h3DC : douta <= 12'hFFB ;
		12'h3DD : douta <= 12'hFFC ;
		12'h3DE : douta <= 12'hFFC ;
		12'h3DF : douta <= 12'hFFC ;
		12'h3E0 : douta <= 12'hFFC ;
		12'h3E1 : douta <= 12'hFFC ;
		12'h3E2 : douta <= 12'hFFC ;
		12'h3E3 : douta <= 12'hFFC ;
		12'h3E4 : douta <= 12'hFFD ;
		12'h3E5 : douta <= 12'hFFD ;
		12'h3E6 : douta <= 12'hFFD ;
		12'h3E7 : douta <= 12'hFFD ;
		12'h3E8 : douta <= 12'hFFD ;
		12'h3E9 : douta <= 12'hFFD ;
		12'h3EA : douta <= 12'hFFD ;
		12'h3EB : douta <= 12'hFFD ;
		12'h3EC : douta <= 12'hFFE ;
		12'h3ED : douta <= 12'hFFE ;
		12'h3EE : douta <= 12'hFFE ;
		12'h3EF : douta <= 12'hFFE ;
		12'h3F0 : douta <= 12'hFFE ;
		12'h3F1 : douta <= 12'hFFE ;
		12'h3F2 : douta <= 12'hFFE ;
		12'h3F3 : douta <= 12'hFFE ;
		12'h3F4 : douta <= 12'hFFE ;
		12'h3F5 : douta <= 12'hFFE ;
		12'h3F6 : douta <= 12'hFFE ;
		12'h3F7 : douta <= 12'hFFE ;
		12'h3F8 : douta <= 12'hFFE ;
		12'h3F9 : douta <= 12'hFFE ;
		12'h3FA : douta <= 12'hFFE ;
		12'h3FB : douta <= 12'hFFE ;
		12'h3FC : douta <= 12'hFFE ;
		12'h3FD : douta <= 12'hFFE ;
		12'h3FE : douta <= 12'hFFE ;
		12'h3FF : douta <= 12'hFFE ;
		12'h400 : douta <= 12'hFFF ;
		12'h401 : douta <= 12'hFFE ;
		12'h402 : douta <= 12'hFFE ;
		12'h403 : douta <= 12'hFFE ;
		12'h404 : douta <= 12'hFFE ;
		12'h405 : douta <= 12'hFFE ;
		12'h406 : douta <= 12'hFFE ;
		12'h407 : douta <= 12'hFFE ;
		12'h408 : douta <= 12'hFFE ;
		12'h409 : douta <= 12'hFFE ;
		12'h40A : douta <= 12'hFFE ;
		12'h40B : douta <= 12'hFFE ;
		12'h40C : douta <= 12'hFFE ;
		12'h40D : douta <= 12'hFFE ;
		12'h40E : douta <= 12'hFFE ;
		12'h40F : douta <= 12'hFFE ;
		12'h410 : douta <= 12'hFFE ;
		12'h411 : douta <= 12'hFFE ;
		12'h412 : douta <= 12'hFFE ;
		12'h413 : douta <= 12'hFFE ;
		12'h414 : douta <= 12'hFFE ;
		12'h415 : douta <= 12'hFFD ;
		12'h416 : douta <= 12'hFFD ;
		12'h417 : douta <= 12'hFFD ;
		12'h418 : douta <= 12'hFFD ;
		12'h419 : douta <= 12'hFFD ;
		12'h41A : douta <= 12'hFFD ;
		12'h41B : douta <= 12'hFFD ;
		12'h41C : douta <= 12'hFFD ;
		12'h41D : douta <= 12'hFFC ;
		12'h41E : douta <= 12'hFFC ;
		12'h41F : douta <= 12'hFFC ;
		12'h420 : douta <= 12'hFFC ;
		12'h421 : douta <= 12'hFFC ;
		12'h422 : douta <= 12'hFFC ;
		12'h423 : douta <= 12'hFFC ;
		12'h424 : douta <= 12'hFFB ;
		12'h425 : douta <= 12'hFFB ;
		12'h426 : douta <= 12'hFFB ;
		12'h427 : douta <= 12'hFFB ;
		12'h428 : douta <= 12'hFFB ;
		12'h429 : douta <= 12'hFFA ;
		12'h42A : douta <= 12'hFFA ;
		12'h42B : douta <= 12'hFFA ;
		12'h42C : douta <= 12'hFFA ;
		12'h42D : douta <= 12'hFFA ;
		12'h42E : douta <= 12'hFF9 ;
		12'h42F : douta <= 12'hFF9 ;
		12'h430 : douta <= 12'hFF9 ;
		12'h431 : douta <= 12'hFF9 ;
		12'h432 : douta <= 12'hFF8 ;
		12'h433 : douta <= 12'hFF8 ;
		12'h434 : douta <= 12'hFF8 ;
		12'h435 : douta <= 12'hFF8 ;
		12'h436 : douta <= 12'hFF7 ;
		12'h437 : douta <= 12'hFF7 ;
		12'h438 : douta <= 12'hFF7 ;
		12'h439 : douta <= 12'hFF7 ;
		12'h43A : douta <= 12'hFF6 ;
		12'h43B : douta <= 12'hFF6 ;
		12'h43C : douta <= 12'hFF6 ;
		12'h43D : douta <= 12'hFF6 ;
		12'h43E : douta <= 12'hFF5 ;
		12'h43F : douta <= 12'hFF5 ;
		12'h440 : douta <= 12'hFF5 ;
		12'h441 : douta <= 12'hFF4 ;
		12'h442 : douta <= 12'hFF4 ;
		12'h443 : douta <= 12'hFF4 ;
		12'h444 : douta <= 12'hFF3 ;
		12'h445 : douta <= 12'hFF3 ;
		12'h446 : douta <= 12'hFF3 ;
		12'h447 : douta <= 12'hFF2 ;
		12'h448 : douta <= 12'hFF2 ;
		12'h449 : douta <= 12'hFF2 ;
		12'h44A : douta <= 12'hFF1 ;
		12'h44B : douta <= 12'hFF1 ;
		12'h44C : douta <= 12'hFF1 ;
		12'h44D : douta <= 12'hFF0 ;
		12'h44E : douta <= 12'hFF0 ;
		12'h44F : douta <= 12'hFEF ;
		12'h450 : douta <= 12'hFEF ;
		12'h451 : douta <= 12'hFEF ;
		12'h452 : douta <= 12'hFEE ;
		12'h453 : douta <= 12'hFEE ;
		12'h454 : douta <= 12'hFEE ;
		12'h455 : douta <= 12'hFED ;
		12'h456 : douta <= 12'hFED ;
		12'h457 : douta <= 12'hFEC ;
		12'h458 : douta <= 12'hFEC ;
		12'h459 : douta <= 12'hFEB ;
		12'h45A : douta <= 12'hFEB ;
		12'h45B : douta <= 12'hFEB ;
		12'h45C : douta <= 12'hFEA ;
		12'h45D : douta <= 12'hFEA ;
		12'h45E : douta <= 12'hFE9 ;
		12'h45F : douta <= 12'hFE9 ;
		12'h460 : douta <= 12'hFE8 ;
		12'h461 : douta <= 12'hFE8 ;
		12'h462 : douta <= 12'hFE7 ;
		12'h463 : douta <= 12'hFE7 ;
		12'h464 : douta <= 12'hFE6 ;
		12'h465 : douta <= 12'hFE6 ;
		12'h466 : douta <= 12'hFE5 ;
		12'h467 : douta <= 12'hFE5 ;
		12'h468 : douta <= 12'hFE5 ;
		12'h469 : douta <= 12'hFE4 ;
		12'h46A : douta <= 12'hFE3 ;
		12'h46B : douta <= 12'hFE3 ;
		12'h46C : douta <= 12'hFE2 ;
		12'h46D : douta <= 12'hFE2 ;
		12'h46E : douta <= 12'hFE1 ;
		12'h46F : douta <= 12'hFE1 ;
		12'h470 : douta <= 12'hFE0 ;
		12'h471 : douta <= 12'hFE0 ;
		12'h472 : douta <= 12'hFDF ;
		12'h473 : douta <= 12'hFDF ;
		12'h474 : douta <= 12'hFDE ;
		12'h475 : douta <= 12'hFDE ;
		12'h476 : douta <= 12'hFDD ;
		12'h477 : douta <= 12'hFDC ;
		12'h478 : douta <= 12'hFDC ;
		12'h479 : douta <= 12'hFDB ;
		12'h47A : douta <= 12'hFDB ;
		12'h47B : douta <= 12'hFDA ;
		12'h47C : douta <= 12'hFDA ;
		12'h47D : douta <= 12'hFD9 ;
		12'h47E : douta <= 12'hFD8 ;
		12'h47F : douta <= 12'hFD8 ;
		12'h480 : douta <= 12'hFD7 ;
		12'h481 : douta <= 12'hFD7 ;
		12'h482 : douta <= 12'hFD6 ;
		12'h483 : douta <= 12'hFD5 ;
		12'h484 : douta <= 12'hFD5 ;
		12'h485 : douta <= 12'hFD4 ;
		12'h486 : douta <= 12'hFD3 ;
		12'h487 : douta <= 12'hFD3 ;
		12'h488 : douta <= 12'hFD2 ;
		12'h489 : douta <= 12'hFD1 ;
		12'h48A : douta <= 12'hFD1 ;
		12'h48B : douta <= 12'hFD0 ;
		12'h48C : douta <= 12'hFCF ;
		12'h48D : douta <= 12'hFCF ;
		12'h48E : douta <= 12'hFCE ;
		12'h48F : douta <= 12'hFCD ;
		12'h490 : douta <= 12'hFCD ;
		12'h491 : douta <= 12'hFCC ;
		12'h492 : douta <= 12'hFCB ;
		12'h493 : douta <= 12'hFCB ;
		12'h494 : douta <= 12'hFCA ;
		12'h495 : douta <= 12'hFC9 ;
		12'h496 : douta <= 12'hFC9 ;
		12'h497 : douta <= 12'hFC8 ;
		12'h498 : douta <= 12'hFC7 ;
		12'h499 : douta <= 12'hFC6 ;
		12'h49A : douta <= 12'hFC6 ;
		12'h49B : douta <= 12'hFC5 ;
		12'h49C : douta <= 12'hFC4 ;
		12'h49D : douta <= 12'hFC3 ;
		12'h49E : douta <= 12'hFC3 ;
		12'h49F : douta <= 12'hFC2 ;
		12'h4A0 : douta <= 12'hFC1 ;
		12'h4A1 : douta <= 12'hFC0 ;
		12'h4A2 : douta <= 12'hFC0 ;
		12'h4A3 : douta <= 12'hFBF ;
		12'h4A4 : douta <= 12'hFBE ;
		12'h4A5 : douta <= 12'hFBD ;
		12'h4A6 : douta <= 12'hFBC ;
		12'h4A7 : douta <= 12'hFBC ;
		12'h4A8 : douta <= 12'hFBB ;
		12'h4A9 : douta <= 12'hFBA ;
		12'h4AA : douta <= 12'hFB9 ;
		12'h4AB : douta <= 12'hFB8 ;
		12'h4AC : douta <= 12'hFB8 ;
		12'h4AD : douta <= 12'hFB7 ;
		12'h4AE : douta <= 12'hFB6 ;
		12'h4AF : douta <= 12'hFB5 ;
		12'h4B0 : douta <= 12'hFB4 ;
		12'h4B1 : douta <= 12'hFB4 ;
		12'h4B2 : douta <= 12'hFB3 ;
		12'h4B3 : douta <= 12'hFB2 ;
		12'h4B4 : douta <= 12'hFB1 ;
		12'h4B5 : douta <= 12'hFB0 ;
		12'h4B6 : douta <= 12'hFAF ;
		12'h4B7 : douta <= 12'hFAE ;
		12'h4B8 : douta <= 12'hFAE ;
		12'h4B9 : douta <= 12'hFAD ;
		12'h4BA : douta <= 12'hFAC ;
		12'h4BB : douta <= 12'hFAB ;
		12'h4BC : douta <= 12'hFAA ;
		12'h4BD : douta <= 12'hFA9 ;
		12'h4BE : douta <= 12'hFA8 ;
		12'h4BF : douta <= 12'hFA7 ;
		12'h4C0 : douta <= 12'hFA6 ;
		12'h4C1 : douta <= 12'hFA5 ;
		12'h4C2 : douta <= 12'hFA5 ;
		12'h4C3 : douta <= 12'hFA4 ;
		12'h4C4 : douta <= 12'hFA3 ;
		12'h4C5 : douta <= 12'hFA2 ;
		12'h4C6 : douta <= 12'hFA1 ;
		12'h4C7 : douta <= 12'hFA0 ;
		12'h4C8 : douta <= 12'hF9F ;
		12'h4C9 : douta <= 12'hF9E ;
		12'h4CA : douta <= 12'hF9D ;
		12'h4CB : douta <= 12'hF9C ;
		12'h4CC : douta <= 12'hF9B ;
		12'h4CD : douta <= 12'hF9A ;
		12'h4CE : douta <= 12'hF99 ;
		12'h4CF : douta <= 12'hF98 ;
		12'h4D0 : douta <= 12'hF97 ;
		12'h4D1 : douta <= 12'hF96 ;
		12'h4D2 : douta <= 12'hF95 ;
		12'h4D3 : douta <= 12'hF94 ;
		12'h4D4 : douta <= 12'hF93 ;
		12'h4D5 : douta <= 12'hF92 ;
		12'h4D6 : douta <= 12'hF91 ;
		12'h4D7 : douta <= 12'hF90 ;
		12'h4D8 : douta <= 12'hF8F ;
		12'h4D9 : douta <= 12'hF8E ;
		12'h4DA : douta <= 12'hF8D ;
		12'h4DB : douta <= 12'hF8C ;
		12'h4DC : douta <= 12'hF8B ;
		12'h4DD : douta <= 12'hF8A ;
		12'h4DE : douta <= 12'hF89 ;
		12'h4DF : douta <= 12'hF88 ;
		12'h4E0 : douta <= 12'hF87 ;
		12'h4E1 : douta <= 12'hF86 ;
		12'h4E2 : douta <= 12'hF85 ;
		12'h4E3 : douta <= 12'hF84 ;
		12'h4E4 : douta <= 12'hF83 ;
		12'h4E5 : douta <= 12'hF81 ;
		12'h4E6 : douta <= 12'hF80 ;
		12'h4E7 : douta <= 12'hF7F ;
		12'h4E8 : douta <= 12'hF7E ;
		12'h4E9 : douta <= 12'hF7D ;
		12'h4EA : douta <= 12'hF7C ;
		12'h4EB : douta <= 12'hF7B ;
		12'h4EC : douta <= 12'hF7A ;
		12'h4ED : douta <= 12'hF79 ;
		12'h4EE : douta <= 12'hF78 ;
		12'h4EF : douta <= 12'hF76 ;
		12'h4F0 : douta <= 12'hF75 ;
		12'h4F1 : douta <= 12'hF74 ;
		12'h4F2 : douta <= 12'hF73 ;
		12'h4F3 : douta <= 12'hF72 ;
		12'h4F4 : douta <= 12'hF71 ;
		12'h4F5 : douta <= 12'hF70 ;
		12'h4F6 : douta <= 12'hF6E ;
		12'h4F7 : douta <= 12'hF6D ;
		12'h4F8 : douta <= 12'hF6C ;
		12'h4F9 : douta <= 12'hF6B ;
		12'h4FA : douta <= 12'hF6A ;
		12'h4FB : douta <= 12'hF69 ;
		12'h4FC : douta <= 12'hF67 ;
		12'h4FD : douta <= 12'hF66 ;
		12'h4FE : douta <= 12'hF65 ;
		12'h4FF : douta <= 12'hF64 ;
		12'h500 : douta <= 12'hF63 ;
		12'h501 : douta <= 12'hF61 ;
		12'h502 : douta <= 12'hF60 ;
		12'h503 : douta <= 12'hF5F ;
		12'h504 : douta <= 12'hF5E ;
		12'h505 : douta <= 12'hF5D ;
		12'h506 : douta <= 12'hF5B ;
		12'h507 : douta <= 12'hF5A ;
		12'h508 : douta <= 12'hF59 ;
		12'h509 : douta <= 12'hF58 ;
		12'h50A : douta <= 12'hF56 ;
		12'h50B : douta <= 12'hF55 ;
		12'h50C : douta <= 12'hF54 ;
		12'h50D : douta <= 12'hF53 ;
		12'h50E : douta <= 12'hF51 ;
		12'h50F : douta <= 12'hF50 ;
		12'h510 : douta <= 12'hF4F ;
		12'h511 : douta <= 12'hF4E ;
		12'h512 : douta <= 12'hF4C ;
		12'h513 : douta <= 12'hF4B ;
		12'h514 : douta <= 12'hF4A ;
		12'h515 : douta <= 12'hF48 ;
		12'h516 : douta <= 12'hF47 ;
		12'h517 : douta <= 12'hF46 ;
		12'h518 : douta <= 12'hF45 ;
		12'h519 : douta <= 12'hF43 ;
		12'h51A : douta <= 12'hF42 ;
		12'h51B : douta <= 12'hF41 ;
		12'h51C : douta <= 12'hF3F ;
		12'h51D : douta <= 12'hF3E ;
		12'h51E : douta <= 12'hF3D ;
		12'h51F : douta <= 12'hF3B ;
		12'h520 : douta <= 12'hF3A ;
		12'h521 : douta <= 12'hF39 ;
		12'h522 : douta <= 12'hF37 ;
		12'h523 : douta <= 12'hF36 ;
		12'h524 : douta <= 12'hF35 ;
		12'h525 : douta <= 12'hF33 ;
		12'h526 : douta <= 12'hF32 ;
		12'h527 : douta <= 12'hF30 ;
		12'h528 : douta <= 12'hF2F ;
		12'h529 : douta <= 12'hF2E ;
		12'h52A : douta <= 12'hF2C ;
		12'h52B : douta <= 12'hF2B ;
		12'h52C : douta <= 12'hF2A ;
		12'h52D : douta <= 12'hF28 ;
		12'h52E : douta <= 12'hF27 ;
		12'h52F : douta <= 12'hF25 ;
		12'h530 : douta <= 12'hF24 ;
		12'h531 : douta <= 12'hF23 ;
		12'h532 : douta <= 12'hF21 ;
		12'h533 : douta <= 12'hF20 ;
		12'h534 : douta <= 12'hF1E ;
		12'h535 : douta <= 12'hF1D ;
		12'h536 : douta <= 12'hF1B ;
		12'h537 : douta <= 12'hF1A ;
		12'h538 : douta <= 12'hF18 ;
		12'h539 : douta <= 12'hF17 ;
		12'h53A : douta <= 12'hF16 ;
		12'h53B : douta <= 12'hF14 ;
		12'h53C : douta <= 12'hF13 ;
		12'h53D : douta <= 12'hF11 ;
		12'h53E : douta <= 12'hF10 ;
		12'h53F : douta <= 12'hF0E ;
		12'h540 : douta <= 12'hF0D ;
		12'h541 : douta <= 12'hF0B ;
		12'h542 : douta <= 12'hF0A ;
		12'h543 : douta <= 12'hF08 ;
		12'h544 : douta <= 12'hF07 ;
		12'h545 : douta <= 12'hF05 ;
		12'h546 : douta <= 12'hF04 ;
		12'h547 : douta <= 12'hF02 ;
		12'h548 : douta <= 12'hF01 ;
		12'h549 : douta <= 12'hEFF ;
		12'h54A : douta <= 12'hEFE ;
		12'h54B : douta <= 12'hEFC ;
		12'h54C : douta <= 12'hEFB ;
		12'h54D : douta <= 12'hEF9 ;
		12'h54E : douta <= 12'hEF8 ;
		12'h54F : douta <= 12'hEF6 ;
		12'h550 : douta <= 12'hEF5 ;
		12'h551 : douta <= 12'hEF3 ;
		12'h552 : douta <= 12'hEF1 ;
		12'h553 : douta <= 12'hEF0 ;
		12'h554 : douta <= 12'hEEE ;
		12'h555 : douta <= 12'hEED ;
		12'h556 : douta <= 12'hEEB ;
		12'h557 : douta <= 12'hEEA ;
		12'h558 : douta <= 12'hEE8 ;
		12'h559 : douta <= 12'hEE6 ;
		12'h55A : douta <= 12'hEE5 ;
		12'h55B : douta <= 12'hEE3 ;
		12'h55C : douta <= 12'hEE2 ;
		12'h55D : douta <= 12'hEE0 ;
		12'h55E : douta <= 12'hEDE ;
		12'h55F : douta <= 12'hEDD ;
		12'h560 : douta <= 12'hEDB ;
		12'h561 : douta <= 12'hEDA ;
		12'h562 : douta <= 12'hED8 ;
		12'h563 : douta <= 12'hED6 ;
		12'h564 : douta <= 12'hED5 ;
		12'h565 : douta <= 12'hED3 ;
		12'h566 : douta <= 12'hED2 ;
		12'h567 : douta <= 12'hED0 ;
		12'h568 : douta <= 12'hECE ;
		12'h569 : douta <= 12'hECD ;
		12'h56A : douta <= 12'hECB ;
		12'h56B : douta <= 12'hEC9 ;
		12'h56C : douta <= 12'hEC8 ;
		12'h56D : douta <= 12'hEC6 ;
		12'h56E : douta <= 12'hEC4 ;
		12'h56F : douta <= 12'hEC3 ;
		12'h570 : douta <= 12'hEC1 ;
		12'h571 : douta <= 12'hEBF ;
		12'h572 : douta <= 12'hEBE ;
		12'h573 : douta <= 12'hEBC ;
		12'h574 : douta <= 12'hEBA ;
		12'h575 : douta <= 12'hEB8 ;
		12'h576 : douta <= 12'hEB7 ;
		12'h577 : douta <= 12'hEB5 ;
		12'h578 : douta <= 12'hEB3 ;
		12'h579 : douta <= 12'hEB2 ;
		12'h57A : douta <= 12'hEB0 ;
		12'h57B : douta <= 12'hEAE ;
		12'h57C : douta <= 12'hEAC ;
		12'h57D : douta <= 12'hEAB ;
		12'h57E : douta <= 12'hEA9 ;
		12'h57F : douta <= 12'hEA7 ;
		12'h580 : douta <= 12'hEA6 ;
		12'h581 : douta <= 12'hEA4 ;
		12'h582 : douta <= 12'hEA2 ;
		12'h583 : douta <= 12'hEA0 ;
		12'h584 : douta <= 12'hE9F ;
		12'h585 : douta <= 12'hE9D ;
		12'h586 : douta <= 12'hE9B ;
		12'h587 : douta <= 12'hE99 ;
		12'h588 : douta <= 12'hE97 ;
		12'h589 : douta <= 12'hE96 ;
		12'h58A : douta <= 12'hE94 ;
		12'h58B : douta <= 12'hE92 ;
		12'h58C : douta <= 12'hE90 ;
		12'h58D : douta <= 12'hE8F ;
		12'h58E : douta <= 12'hE8D ;
		12'h58F : douta <= 12'hE8B ;
		12'h590 : douta <= 12'hE89 ;
		12'h591 : douta <= 12'hE87 ;
		12'h592 : douta <= 12'hE85 ;
		12'h593 : douta <= 12'hE84 ;
		12'h594 : douta <= 12'hE82 ;
		12'h595 : douta <= 12'hE80 ;
		12'h596 : douta <= 12'hE7E ;
		12'h597 : douta <= 12'hE7C ;
		12'h598 : douta <= 12'hE7B ;
		12'h599 : douta <= 12'hE79 ;
		12'h59A : douta <= 12'hE77 ;
		12'h59B : douta <= 12'hE75 ;
		12'h59C : douta <= 12'hE73 ;
		12'h59D : douta <= 12'hE71 ;
		12'h59E : douta <= 12'hE6F ;
		12'h59F : douta <= 12'hE6E ;
		12'h5A0 : douta <= 12'hE6C ;
		12'h5A1 : douta <= 12'hE6A ;
		12'h5A2 : douta <= 12'hE68 ;
		12'h5A3 : douta <= 12'hE66 ;
		12'h5A4 : douta <= 12'hE64 ;
		12'h5A5 : douta <= 12'hE62 ;
		12'h5A6 : douta <= 12'hE60 ;
		12'h5A7 : douta <= 12'hE5E ;
		12'h5A8 : douta <= 12'hE5D ;
		12'h5A9 : douta <= 12'hE5B ;
		12'h5AA : douta <= 12'hE59 ;
		12'h5AB : douta <= 12'hE57 ;
		12'h5AC : douta <= 12'hE55 ;
		12'h5AD : douta <= 12'hE53 ;
		12'h5AE : douta <= 12'hE51 ;
		12'h5AF : douta <= 12'hE4F ;
		12'h5B0 : douta <= 12'hE4D ;
		12'h5B1 : douta <= 12'hE4B ;
		12'h5B2 : douta <= 12'hE49 ;
		12'h5B3 : douta <= 12'hE47 ;
		12'h5B4 : douta <= 12'hE45 ;
		12'h5B5 : douta <= 12'hE44 ;
		12'h5B6 : douta <= 12'hE42 ;
		12'h5B7 : douta <= 12'hE40 ;
		12'h5B8 : douta <= 12'hE3E ;
		12'h5B9 : douta <= 12'hE3C ;
		12'h5BA : douta <= 12'hE3A ;
		12'h5BB : douta <= 12'hE38 ;
		12'h5BC : douta <= 12'hE36 ;
		12'h5BD : douta <= 12'hE34 ;
		12'h5BE : douta <= 12'hE32 ;
		12'h5BF : douta <= 12'hE30 ;
		12'h5C0 : douta <= 12'hE2E ;
		12'h5C1 : douta <= 12'hE2C ;
		12'h5C2 : douta <= 12'hE2A ;
		12'h5C3 : douta <= 12'hE28 ;
		12'h5C4 : douta <= 12'hE26 ;
		12'h5C5 : douta <= 12'hE24 ;
		12'h5C6 : douta <= 12'hE22 ;
		12'h5C7 : douta <= 12'hE20 ;
		12'h5C8 : douta <= 12'hE1E ;
		12'h5C9 : douta <= 12'hE1C ;
		12'h5CA : douta <= 12'hE1A ;
		12'h5CB : douta <= 12'hE18 ;
		12'h5CC : douta <= 12'hE16 ;
		12'h5CD : douta <= 12'hE14 ;
		12'h5CE : douta <= 12'hE12 ;
		12'h5CF : douta <= 12'hE10 ;
		12'h5D0 : douta <= 12'hE0E ;
		12'h5D1 : douta <= 12'hE0B ;
		12'h5D2 : douta <= 12'hE09 ;
		12'h5D3 : douta <= 12'hE07 ;
		12'h5D4 : douta <= 12'hE05 ;
		12'h5D5 : douta <= 12'hE03 ;
		12'h5D6 : douta <= 12'hE01 ;
		12'h5D7 : douta <= 12'hDFF ;
		12'h5D8 : douta <= 12'hDFD ;
		12'h5D9 : douta <= 12'hDFB ;
		12'h5DA : douta <= 12'hDF9 ;
		12'h5DB : douta <= 12'hDF7 ;
		12'h5DC : douta <= 12'hDF5 ;
		12'h5DD : douta <= 12'hDF3 ;
		12'h5DE : douta <= 12'hDF0 ;
		12'h5DF : douta <= 12'hDEE ;
		12'h5E0 : douta <= 12'hDEC ;
		12'h5E1 : douta <= 12'hDEA ;
		12'h5E2 : douta <= 12'hDE8 ;
		12'h5E3 : douta <= 12'hDE6 ;
		12'h5E4 : douta <= 12'hDE4 ;
		12'h5E5 : douta <= 12'hDE2 ;
		12'h5E6 : douta <= 12'hDE0 ;
		12'h5E7 : douta <= 12'hDDD ;
		12'h5E8 : douta <= 12'hDDB ;
		12'h5E9 : douta <= 12'hDD9 ;
		12'h5EA : douta <= 12'hDD7 ;
		12'h5EB : douta <= 12'hDD5 ;
		12'h5EC : douta <= 12'hDD3 ;
		12'h5ED : douta <= 12'hDD1 ;
		12'h5EE : douta <= 12'hDCE ;
		12'h5EF : douta <= 12'hDCC ;
		12'h5F0 : douta <= 12'hDCA ;
		12'h5F1 : douta <= 12'hDC8 ;
		12'h5F2 : douta <= 12'hDC6 ;
		12'h5F3 : douta <= 12'hDC4 ;
		12'h5F4 : douta <= 12'hDC1 ;
		12'h5F5 : douta <= 12'hDBF ;
		12'h5F6 : douta <= 12'hDBD ;
		12'h5F7 : douta <= 12'hDBB ;
		12'h5F8 : douta <= 12'hDB9 ;
		12'h5F9 : douta <= 12'hDB6 ;
		12'h5FA : douta <= 12'hDB4 ;
		12'h5FB : douta <= 12'hDB2 ;
		12'h5FC : douta <= 12'hDB0 ;
		12'h5FD : douta <= 12'hDAE ;
		12'h5FE : douta <= 12'hDAB ;
		12'h5FF : douta <= 12'hDA9 ;
		12'h600 : douta <= 12'hDA7 ;
		12'h601 : douta <= 12'hDA5 ;
		12'h602 : douta <= 12'hDA3 ;
		12'h603 : douta <= 12'hDA0 ;
		12'h604 : douta <= 12'hD9E ;
		12'h605 : douta <= 12'hD9C ;
		12'h606 : douta <= 12'hD9A ;
		12'h607 : douta <= 12'hD97 ;
		12'h608 : douta <= 12'hD95 ;
		12'h609 : douta <= 12'hD93 ;
		12'h60A : douta <= 12'hD91 ;
		12'h60B : douta <= 12'hD8E ;
		12'h60C : douta <= 12'hD8C ;
		12'h60D : douta <= 12'hD8A ;
		12'h60E : douta <= 12'hD88 ;
		12'h60F : douta <= 12'hD85 ;
		12'h610 : douta <= 12'hD83 ;
		12'h611 : douta <= 12'hD81 ;
		12'h612 : douta <= 12'hD7E ;
		12'h613 : douta <= 12'hD7C ;
		12'h614 : douta <= 12'hD7A ;
		12'h615 : douta <= 12'hD78 ;
		12'h616 : douta <= 12'hD75 ;
		12'h617 : douta <= 12'hD73 ;
		12'h618 : douta <= 12'hD71 ;
		12'h619 : douta <= 12'hD6E ;
		12'h61A : douta <= 12'hD6C ;
		12'h61B : douta <= 12'hD6A ;
		12'h61C : douta <= 12'hD67 ;
		12'h61D : douta <= 12'hD65 ;
		12'h61E : douta <= 12'hD63 ;
		12'h61F : douta <= 12'hD61 ;
		12'h620 : douta <= 12'hD5E ;
		12'h621 : douta <= 12'hD5C ;
		12'h622 : douta <= 12'hD5A ;
		12'h623 : douta <= 12'hD57 ;
		12'h624 : douta <= 12'hD55 ;
		12'h625 : douta <= 12'hD53 ;
		12'h626 : douta <= 12'hD50 ;
		12'h627 : douta <= 12'hD4E ;
		12'h628 : douta <= 12'hD4B ;
		12'h629 : douta <= 12'hD49 ;
		12'h62A : douta <= 12'hD47 ;
		12'h62B : douta <= 12'hD44 ;
		12'h62C : douta <= 12'hD42 ;
		12'h62D : douta <= 12'hD40 ;
		12'h62E : douta <= 12'hD3D ;
		12'h62F : douta <= 12'hD3B ;
		12'h630 : douta <= 12'hD39 ;
		12'h631 : douta <= 12'hD36 ;
		12'h632 : douta <= 12'hD34 ;
		12'h633 : douta <= 12'hD31 ;
		12'h634 : douta <= 12'hD2F ;
		12'h635 : douta <= 12'hD2D ;
		12'h636 : douta <= 12'hD2A ;
		12'h637 : douta <= 12'hD28 ;
		12'h638 : douta <= 12'hD25 ;
		12'h639 : douta <= 12'hD23 ;
		12'h63A : douta <= 12'hD21 ;
		12'h63B : douta <= 12'hD1E ;
		12'h63C : douta <= 12'hD1C ;
		12'h63D : douta <= 12'hD19 ;
		12'h63E : douta <= 12'hD17 ;
		12'h63F : douta <= 12'hD15 ;
		12'h640 : douta <= 12'hD12 ;
		12'h641 : douta <= 12'hD10 ;
		12'h642 : douta <= 12'hD0D ;
		12'h643 : douta <= 12'hD0B ;
		12'h644 : douta <= 12'hD08 ;
		12'h645 : douta <= 12'hD06 ;
		12'h646 : douta <= 12'hD03 ;
		12'h647 : douta <= 12'hD01 ;
		12'h648 : douta <= 12'hCFF ;
		12'h649 : douta <= 12'hCFC ;
		12'h64A : douta <= 12'hCFA ;
		12'h64B : douta <= 12'hCF7 ;
		12'h64C : douta <= 12'hCF5 ;
		12'h64D : douta <= 12'hCF2 ;
		12'h64E : douta <= 12'hCF0 ;
		12'h64F : douta <= 12'hCED ;
		12'h650 : douta <= 12'hCEB ;
		12'h651 : douta <= 12'hCE8 ;
		12'h652 : douta <= 12'hCE6 ;
		12'h653 : douta <= 12'hCE3 ;
		12'h654 : douta <= 12'hCE1 ;
		12'h655 : douta <= 12'hCDE ;
		12'h656 : douta <= 12'hCDC ;
		12'h657 : douta <= 12'hCD9 ;
		12'h658 : douta <= 12'hCD7 ;
		12'h659 : douta <= 12'hCD4 ;
		12'h65A : douta <= 12'hCD2 ;
		12'h65B : douta <= 12'hCCF ;
		12'h65C : douta <= 12'hCCD ;
		12'h65D : douta <= 12'hCCA ;
		12'h65E : douta <= 12'hCC8 ;
		12'h65F : douta <= 12'hCC5 ;
		12'h660 : douta <= 12'hCC3 ;
		12'h661 : douta <= 12'hCC0 ;
		12'h662 : douta <= 12'hCBE ;
		12'h663 : douta <= 12'hCBB ;
		12'h664 : douta <= 12'hCB9 ;
		12'h665 : douta <= 12'hCB6 ;
		12'h666 : douta <= 12'hCB4 ;
		12'h667 : douta <= 12'hCB1 ;
		12'h668 : douta <= 12'hCAF ;
		12'h669 : douta <= 12'hCAC ;
		12'h66A : douta <= 12'hCAA ;
		12'h66B : douta <= 12'hCA7 ;
		12'h66C : douta <= 12'hCA4 ;
		12'h66D : douta <= 12'hCA2 ;
		12'h66E : douta <= 12'hC9F ;
		12'h66F : douta <= 12'hC9D ;
		12'h670 : douta <= 12'hC9A ;
		12'h671 : douta <= 12'hC98 ;
		12'h672 : douta <= 12'hC95 ;
		12'h673 : douta <= 12'hC92 ;
		12'h674 : douta <= 12'hC90 ;
		12'h675 : douta <= 12'hC8D ;
		12'h676 : douta <= 12'hC8B ;
		12'h677 : douta <= 12'hC88 ;
		12'h678 : douta <= 12'hC86 ;
		12'h679 : douta <= 12'hC83 ;
		12'h67A : douta <= 12'hC80 ;
		12'h67B : douta <= 12'hC7E ;
		12'h67C : douta <= 12'hC7B ;
		12'h67D : douta <= 12'hC79 ;
		12'h67E : douta <= 12'hC76 ;
		12'h67F : douta <= 12'hC73 ;
		12'h680 : douta <= 12'hC71 ;
		12'h681 : douta <= 12'hC6E ;
		12'h682 : douta <= 12'hC6C ;
		12'h683 : douta <= 12'hC69 ;
		12'h684 : douta <= 12'hC66 ;
		12'h685 : douta <= 12'hC64 ;
		12'h686 : douta <= 12'hC61 ;
		12'h687 : douta <= 12'hC5E ;
		12'h688 : douta <= 12'hC5C ;
		12'h689 : douta <= 12'hC59 ;
		12'h68A : douta <= 12'hC57 ;
		12'h68B : douta <= 12'hC54 ;
		12'h68C : douta <= 12'hC51 ;
		12'h68D : douta <= 12'hC4F ;
		12'h68E : douta <= 12'hC4C ;
		12'h68F : douta <= 12'hC49 ;
		12'h690 : douta <= 12'hC47 ;
		12'h691 : douta <= 12'hC44 ;
		12'h692 : douta <= 12'hC41 ;
		12'h693 : douta <= 12'hC3F ;
		12'h694 : douta <= 12'hC3C ;
		12'h695 : douta <= 12'hC39 ;
		12'h696 : douta <= 12'hC37 ;
		12'h697 : douta <= 12'hC34 ;
		12'h698 : douta <= 12'hC31 ;
		12'h699 : douta <= 12'hC2F ;
		12'h69A : douta <= 12'hC2C ;
		12'h69B : douta <= 12'hC29 ;
		12'h69C : douta <= 12'hC27 ;
		12'h69D : douta <= 12'hC24 ;
		12'h69E : douta <= 12'hC21 ;
		12'h69F : douta <= 12'hC1F ;
		12'h6A0 : douta <= 12'hC1C ;
		12'h6A1 : douta <= 12'hC19 ;
		12'h6A2 : douta <= 12'hC16 ;
		12'h6A3 : douta <= 12'hC14 ;
		12'h6A4 : douta <= 12'hC11 ;
		12'h6A5 : douta <= 12'hC0E ;
		12'h6A6 : douta <= 12'hC0C ;
		12'h6A7 : douta <= 12'hC09 ;
		12'h6A8 : douta <= 12'hC06 ;
		12'h6A9 : douta <= 12'hC04 ;
		12'h6AA : douta <= 12'hC01 ;
		12'h6AB : douta <= 12'hBFE ;
		12'h6AC : douta <= 12'hBFB ;
		12'h6AD : douta <= 12'hBF9 ;
		12'h6AE : douta <= 12'hBF6 ;
		12'h6AF : douta <= 12'hBF3 ;
		12'h6B0 : douta <= 12'hBF0 ;
		12'h6B1 : douta <= 12'hBEE ;
		12'h6B2 : douta <= 12'hBEB ;
		12'h6B3 : douta <= 12'hBE8 ;
		12'h6B4 : douta <= 12'hBE6 ;
		12'h6B5 : douta <= 12'hBE3 ;
		12'h6B6 : douta <= 12'hBE0 ;
		12'h6B7 : douta <= 12'hBDD ;
		12'h6B8 : douta <= 12'hBDB ;
		12'h6B9 : douta <= 12'hBD8 ;
		12'h6BA : douta <= 12'hBD5 ;
		12'h6BB : douta <= 12'hBD2 ;
		12'h6BC : douta <= 12'hBD0 ;
		12'h6BD : douta <= 12'hBCD ;
		12'h6BE : douta <= 12'hBCA ;
		12'h6BF : douta <= 12'hBC7 ;
		12'h6C0 : douta <= 12'hBC4 ;
		12'h6C1 : douta <= 12'hBC2 ;
		12'h6C2 : douta <= 12'hBBF ;
		12'h6C3 : douta <= 12'hBBC ;
		12'h6C4 : douta <= 12'hBB9 ;
		12'h6C5 : douta <= 12'hBB7 ;
		12'h6C6 : douta <= 12'hBB4 ;
		12'h6C7 : douta <= 12'hBB1 ;
		12'h6C8 : douta <= 12'hBAE ;
		12'h6C9 : douta <= 12'hBAB ;
		12'h6CA : douta <= 12'hBA9 ;
		12'h6CB : douta <= 12'hBA6 ;
		12'h6CC : douta <= 12'hBA3 ;
		12'h6CD : douta <= 12'hBA0 ;
		12'h6CE : douta <= 12'hB9D ;
		12'h6CF : douta <= 12'hB9B ;
		12'h6D0 : douta <= 12'hB98 ;
		12'h6D1 : douta <= 12'hB95 ;
		12'h6D2 : douta <= 12'hB92 ;
		12'h6D3 : douta <= 12'hB8F ;
		12'h6D4 : douta <= 12'hB8D ;
		12'h6D5 : douta <= 12'hB8A ;
		12'h6D6 : douta <= 12'hB87 ;
		12'h6D7 : douta <= 12'hB84 ;
		12'h6D8 : douta <= 12'hB81 ;
		12'h6D9 : douta <= 12'hB7F ;
		12'h6DA : douta <= 12'hB7C ;
		12'h6DB : douta <= 12'hB79 ;
		12'h6DC : douta <= 12'hB76 ;
		12'h6DD : douta <= 12'hB73 ;
		12'h6DE : douta <= 12'hB70 ;
		12'h6DF : douta <= 12'hB6E ;
		12'h6E0 : douta <= 12'hB6B ;
		12'h6E1 : douta <= 12'hB68 ;
		12'h6E2 : douta <= 12'hB65 ;
		12'h6E3 : douta <= 12'hB62 ;
		12'h6E4 : douta <= 12'hB5F ;
		12'h6E5 : douta <= 12'hB5C ;
		12'h6E6 : douta <= 12'hB5A ;
		12'h6E7 : douta <= 12'hB57 ;
		12'h6E8 : douta <= 12'hB54 ;
		12'h6E9 : douta <= 12'hB51 ;
		12'h6EA : douta <= 12'hB4E ;
		12'h6EB : douta <= 12'hB4B ;
		12'h6EC : douta <= 12'hB48 ;
		12'h6ED : douta <= 12'hB46 ;
		12'h6EE : douta <= 12'hB43 ;
		12'h6EF : douta <= 12'hB40 ;
		12'h6F0 : douta <= 12'hB3D ;
		12'h6F1 : douta <= 12'hB3A ;
		12'h6F2 : douta <= 12'hB37 ;
		12'h6F3 : douta <= 12'hB34 ;
		12'h6F4 : douta <= 12'hB32 ;
		12'h6F5 : douta <= 12'hB2F ;
		12'h6F6 : douta <= 12'hB2C ;
		12'h6F7 : douta <= 12'hB29 ;
		12'h6F8 : douta <= 12'hB26 ;
		12'h6F9 : douta <= 12'hB23 ;
		12'h6FA : douta <= 12'hB20 ;
		12'h6FB : douta <= 12'hB1D ;
		12'h6FC : douta <= 12'hB1A ;
		12'h6FD : douta <= 12'hB18 ;
		12'h6FE : douta <= 12'hB15 ;
		12'h6FF : douta <= 12'hB12 ;
		12'h700 : douta <= 12'hB0F ;
		12'h701 : douta <= 12'hB0C ;
		12'h702 : douta <= 12'hB09 ;
		12'h703 : douta <= 12'hB06 ;
		12'h704 : douta <= 12'hB03 ;
		12'h705 : douta <= 12'hB00 ;
		12'h706 : douta <= 12'hAFD ;
		12'h707 : douta <= 12'hAFB ;
		12'h708 : douta <= 12'hAF8 ;
		12'h709 : douta <= 12'hAF5 ;
		12'h70A : douta <= 12'hAF2 ;
		12'h70B : douta <= 12'hAEF ;
		12'h70C : douta <= 12'hAEC ;
		12'h70D : douta <= 12'hAE9 ;
		12'h70E : douta <= 12'hAE6 ;
		12'h70F : douta <= 12'hAE3 ;
		12'h710 : douta <= 12'hAE0 ;
		12'h711 : douta <= 12'hADD ;
		12'h712 : douta <= 12'hADA ;
		12'h713 : douta <= 12'hAD7 ;
		12'h714 : douta <= 12'hAD4 ;
		12'h715 : douta <= 12'hAD2 ;
		12'h716 : douta <= 12'hACF ;
		12'h717 : douta <= 12'hACC ;
		12'h718 : douta <= 12'hAC9 ;
		12'h719 : douta <= 12'hAC6 ;
		12'h71A : douta <= 12'hAC3 ;
		12'h71B : douta <= 12'hAC0 ;
		12'h71C : douta <= 12'hABD ;
		12'h71D : douta <= 12'hABA ;
		12'h71E : douta <= 12'hAB7 ;
		12'h71F : douta <= 12'hAB4 ;
		12'h720 : douta <= 12'hAB1 ;
		12'h721 : douta <= 12'hAAE ;
		12'h722 : douta <= 12'hAAB ;
		12'h723 : douta <= 12'hAA8 ;
		12'h724 : douta <= 12'hAA5 ;
		12'h725 : douta <= 12'hAA2 ;
		12'h726 : douta <= 12'hA9F ;
		12'h727 : douta <= 12'hA9C ;
		12'h728 : douta <= 12'hA99 ;
		12'h729 : douta <= 12'hA96 ;
		12'h72A : douta <= 12'hA93 ;
		12'h72B : douta <= 12'hA90 ;
		12'h72C : douta <= 12'hA8E ;
		12'h72D : douta <= 12'hA8B ;
		12'h72E : douta <= 12'hA88 ;
		12'h72F : douta <= 12'hA85 ;
		12'h730 : douta <= 12'hA82 ;
		12'h731 : douta <= 12'hA7F ;
		12'h732 : douta <= 12'hA7C ;
		12'h733 : douta <= 12'hA79 ;
		12'h734 : douta <= 12'hA76 ;
		12'h735 : douta <= 12'hA73 ;
		12'h736 : douta <= 12'hA70 ;
		12'h737 : douta <= 12'hA6D ;
		12'h738 : douta <= 12'hA6A ;
		12'h739 : douta <= 12'hA67 ;
		12'h73A : douta <= 12'hA64 ;
		12'h73B : douta <= 12'hA61 ;
		12'h73C : douta <= 12'hA5E ;
		12'h73D : douta <= 12'hA5B ;
		12'h73E : douta <= 12'hA58 ;
		12'h73F : douta <= 12'hA55 ;
		12'h740 : douta <= 12'hA52 ;
		12'h741 : douta <= 12'hA4F ;
		12'h742 : douta <= 12'hA4C ;
		12'h743 : douta <= 12'hA49 ;
		12'h744 : douta <= 12'hA46 ;
		12'h745 : douta <= 12'hA43 ;
		12'h746 : douta <= 12'hA40 ;
		12'h747 : douta <= 12'hA3D ;
		12'h748 : douta <= 12'hA3A ;
		12'h749 : douta <= 12'hA37 ;
		12'h74A : douta <= 12'hA34 ;
		12'h74B : douta <= 12'hA31 ;
		12'h74C : douta <= 12'hA2E ;
		12'h74D : douta <= 12'hA2B ;
		12'h74E : douta <= 12'hA28 ;
		12'h74F : douta <= 12'hA24 ;
		12'h750 : douta <= 12'hA21 ;
		12'h751 : douta <= 12'hA1E ;
		12'h752 : douta <= 12'hA1B ;
		12'h753 : douta <= 12'hA18 ;
		12'h754 : douta <= 12'hA15 ;
		12'h755 : douta <= 12'hA12 ;
		12'h756 : douta <= 12'hA0F ;
		12'h757 : douta <= 12'hA0C ;
		12'h758 : douta <= 12'hA09 ;
		12'h759 : douta <= 12'hA06 ;
		12'h75A : douta <= 12'hA03 ;
		12'h75B : douta <= 12'hA00 ;
		12'h75C : douta <= 12'h9FD ;
		12'h75D : douta <= 12'h9FA ;
		12'h75E : douta <= 12'h9F7 ;
		12'h75F : douta <= 12'h9F4 ;
		12'h760 : douta <= 12'h9F1 ;
		12'h761 : douta <= 12'h9EE ;
		12'h762 : douta <= 12'h9EB ;
		12'h763 : douta <= 12'h9E8 ;
		12'h764 : douta <= 12'h9E5 ;
		12'h765 : douta <= 12'h9E2 ;
		12'h766 : douta <= 12'h9DF ;
		12'h767 : douta <= 12'h9DC ;
		12'h768 : douta <= 12'h9D8 ;
		12'h769 : douta <= 12'h9D5 ;
		12'h76A : douta <= 12'h9D2 ;
		12'h76B : douta <= 12'h9CF ;
		12'h76C : douta <= 12'h9CC ;
		12'h76D : douta <= 12'h9C9 ;
		12'h76E : douta <= 12'h9C6 ;
		12'h76F : douta <= 12'h9C3 ;
		12'h770 : douta <= 12'h9C0 ;
		12'h771 : douta <= 12'h9BD ;
		12'h772 : douta <= 12'h9BA ;
		12'h773 : douta <= 12'h9B7 ;
		12'h774 : douta <= 12'h9B4 ;
		12'h775 : douta <= 12'h9B1 ;
		12'h776 : douta <= 12'h9AE ;
		12'h777 : douta <= 12'h9AB ;
		12'h778 : douta <= 12'h9A7 ;
		12'h779 : douta <= 12'h9A4 ;
		12'h77A : douta <= 12'h9A1 ;
		12'h77B : douta <= 12'h99E ;
		12'h77C : douta <= 12'h99B ;
		12'h77D : douta <= 12'h998 ;
		12'h77E : douta <= 12'h995 ;
		12'h77F : douta <= 12'h992 ;
		12'h780 : douta <= 12'h98F ;
		12'h781 : douta <= 12'h98C ;
		12'h782 : douta <= 12'h989 ;
		12'h783 : douta <= 12'h986 ;
		12'h784 : douta <= 12'h983 ;
		12'h785 : douta <= 12'h97F ;
		12'h786 : douta <= 12'h97C ;
		12'h787 : douta <= 12'h979 ;
		12'h788 : douta <= 12'h976 ;
		12'h789 : douta <= 12'h973 ;
		12'h78A : douta <= 12'h970 ;
		12'h78B : douta <= 12'h96D ;
		12'h78C : douta <= 12'h96A ;
		12'h78D : douta <= 12'h967 ;
		12'h78E : douta <= 12'h964 ;
		12'h78F : douta <= 12'h961 ;
		12'h790 : douta <= 12'h95D ;
		12'h791 : douta <= 12'h95A ;
		12'h792 : douta <= 12'h957 ;
		12'h793 : douta <= 12'h954 ;
		12'h794 : douta <= 12'h951 ;
		12'h795 : douta <= 12'h94E ;
		12'h796 : douta <= 12'h94B ;
		12'h797 : douta <= 12'h948 ;
		12'h798 : douta <= 12'h945 ;
		12'h799 : douta <= 12'h942 ;
		12'h79A : douta <= 12'h93E ;
		12'h79B : douta <= 12'h93B ;
		12'h79C : douta <= 12'h938 ;
		12'h79D : douta <= 12'h935 ;
		12'h79E : douta <= 12'h932 ;
		12'h79F : douta <= 12'h92F ;
		12'h7A0 : douta <= 12'h92C ;
		12'h7A1 : douta <= 12'h929 ;
		12'h7A2 : douta <= 12'h926 ;
		12'h7A3 : douta <= 12'h923 ;
		12'h7A4 : douta <= 12'h91F ;
		12'h7A5 : douta <= 12'h91C ;
		12'h7A6 : douta <= 12'h919 ;
		12'h7A7 : douta <= 12'h916 ;
		12'h7A8 : douta <= 12'h913 ;
		12'h7A9 : douta <= 12'h910 ;
		12'h7AA : douta <= 12'h90D ;
		12'h7AB : douta <= 12'h90A ;
		12'h7AC : douta <= 12'h907 ;
		12'h7AD : douta <= 12'h903 ;
		12'h7AE : douta <= 12'h900 ;
		12'h7AF : douta <= 12'h8FD ;
		12'h7B0 : douta <= 12'h8FA ;
		12'h7B1 : douta <= 12'h8F7 ;
		12'h7B2 : douta <= 12'h8F4 ;
		12'h7B3 : douta <= 12'h8F1 ;
		12'h7B4 : douta <= 12'h8EE ;
		12'h7B5 : douta <= 12'h8EA ;
		12'h7B6 : douta <= 12'h8E7 ;
		12'h7B7 : douta <= 12'h8E4 ;
		12'h7B8 : douta <= 12'h8E1 ;
		12'h7B9 : douta <= 12'h8DE ;
		12'h7BA : douta <= 12'h8DB ;
		12'h7BB : douta <= 12'h8D8 ;
		12'h7BC : douta <= 12'h8D5 ;
		12'h7BD : douta <= 12'h8D2 ;
		12'h7BE : douta <= 12'h8CE ;
		12'h7BF : douta <= 12'h8CB ;
		12'h7C0 : douta <= 12'h8C8 ;
		12'h7C1 : douta <= 12'h8C5 ;
		12'h7C2 : douta <= 12'h8C2 ;
		12'h7C3 : douta <= 12'h8BF ;
		12'h7C4 : douta <= 12'h8BC ;
		12'h7C5 : douta <= 12'h8B9 ;
		12'h7C6 : douta <= 12'h8B5 ;
		12'h7C7 : douta <= 12'h8B2 ;
		12'h7C8 : douta <= 12'h8AF ;
		12'h7C9 : douta <= 12'h8AC ;
		12'h7CA : douta <= 12'h8A9 ;
		12'h7CB : douta <= 12'h8A6 ;
		12'h7CC : douta <= 12'h8A3 ;
		12'h7CD : douta <= 12'h89F ;
		12'h7CE : douta <= 12'h89C ;
		12'h7CF : douta <= 12'h899 ;
		12'h7D0 : douta <= 12'h896 ;
		12'h7D1 : douta <= 12'h893 ;
		12'h7D2 : douta <= 12'h890 ;
		12'h7D3 : douta <= 12'h88D ;
		12'h7D4 : douta <= 12'h88A ;
		12'h7D5 : douta <= 12'h886 ;
		12'h7D6 : douta <= 12'h883 ;
		12'h7D7 : douta <= 12'h880 ;
		12'h7D8 : douta <= 12'h87D ;
		12'h7D9 : douta <= 12'h87A ;
		12'h7DA : douta <= 12'h877 ;
		12'h7DB : douta <= 12'h874 ;
		12'h7DC : douta <= 12'h870 ;
		12'h7DD : douta <= 12'h86D ;
		12'h7DE : douta <= 12'h86A ;
		12'h7DF : douta <= 12'h867 ;
		12'h7E0 : douta <= 12'h864 ;
		12'h7E1 : douta <= 12'h861 ;
		12'h7E2 : douta <= 12'h85E ;
		12'h7E3 : douta <= 12'h85B ;
		12'h7E4 : douta <= 12'h857 ;
		12'h7E5 : douta <= 12'h854 ;
		12'h7E6 : douta <= 12'h851 ;
		12'h7E7 : douta <= 12'h84E ;
		12'h7E8 : douta <= 12'h84B ;
		12'h7E9 : douta <= 12'h848 ;
		12'h7EA : douta <= 12'h845 ;
		12'h7EB : douta <= 12'h841 ;
		12'h7EC : douta <= 12'h83E ;
		12'h7ED : douta <= 12'h83B ;
		12'h7EE : douta <= 12'h838 ;
		12'h7EF : douta <= 12'h835 ;
		12'h7F0 : douta <= 12'h832 ;
		12'h7F1 : douta <= 12'h82F ;
		12'h7F2 : douta <= 12'h82B ;
		12'h7F3 : douta <= 12'h828 ;
		12'h7F4 : douta <= 12'h825 ;
		12'h7F5 : douta <= 12'h822 ;
		12'h7F6 : douta <= 12'h81F ;
		12'h7F7 : douta <= 12'h81C ;
		12'h7F8 : douta <= 12'h819 ;
		12'h7F9 : douta <= 12'h815 ;
		12'h7FA : douta <= 12'h812 ;
		12'h7FB : douta <= 12'h80F ;
		12'h7FC : douta <= 12'h80C ;
		12'h7FD : douta <= 12'h809 ;
		12'h7FE : douta <= 12'h806 ;
		12'h7FF : douta <= 12'h803 ;
		12'h800 : douta <= 12'h800 ;
		12'h801 : douta <= 12'h7FC ;
		12'h802 : douta <= 12'h7F9 ;
		12'h803 : douta <= 12'h7F6 ;
		12'h804 : douta <= 12'h7F3 ;
		12'h805 : douta <= 12'h7F0 ;
		12'h806 : douta <= 12'h7ED ;
		12'h807 : douta <= 12'h7EA ;
		12'h808 : douta <= 12'h7E6 ;
		12'h809 : douta <= 12'h7E3 ;
		12'h80A : douta <= 12'h7E0 ;
		12'h80B : douta <= 12'h7DD ;
		12'h80C : douta <= 12'h7DA ;
		12'h80D : douta <= 12'h7D7 ;
		12'h80E : douta <= 12'h7D4 ;
		12'h80F : douta <= 12'h7D0 ;
		12'h810 : douta <= 12'h7CD ;
		12'h811 : douta <= 12'h7CA ;
		12'h812 : douta <= 12'h7C7 ;
		12'h813 : douta <= 12'h7C4 ;
		12'h814 : douta <= 12'h7C1 ;
		12'h815 : douta <= 12'h7BE ;
		12'h816 : douta <= 12'h7BA ;
		12'h817 : douta <= 12'h7B7 ;
		12'h818 : douta <= 12'h7B4 ;
		12'h819 : douta <= 12'h7B1 ;
		12'h81A : douta <= 12'h7AE ;
		12'h81B : douta <= 12'h7AB ;
		12'h81C : douta <= 12'h7A8 ;
		12'h81D : douta <= 12'h7A4 ;
		12'h81E : douta <= 12'h7A1 ;
		12'h81F : douta <= 12'h79E ;
		12'h820 : douta <= 12'h79B ;
		12'h821 : douta <= 12'h798 ;
		12'h822 : douta <= 12'h795 ;
		12'h823 : douta <= 12'h792 ;
		12'h824 : douta <= 12'h78F ;
		12'h825 : douta <= 12'h78B ;
		12'h826 : douta <= 12'h788 ;
		12'h827 : douta <= 12'h785 ;
		12'h828 : douta <= 12'h782 ;
		12'h829 : douta <= 12'h77F ;
		12'h82A : douta <= 12'h77C ;
		12'h82B : douta <= 12'h779 ;
		12'h82C : douta <= 12'h775 ;
		12'h82D : douta <= 12'h772 ;
		12'h82E : douta <= 12'h76F ;
		12'h82F : douta <= 12'h76C ;
		12'h830 : douta <= 12'h769 ;
		12'h831 : douta <= 12'h766 ;
		12'h832 : douta <= 12'h763 ;
		12'h833 : douta <= 12'h760 ;
		12'h834 : douta <= 12'h75C ;
		12'h835 : douta <= 12'h759 ;
		12'h836 : douta <= 12'h756 ;
		12'h837 : douta <= 12'h753 ;
		12'h838 : douta <= 12'h750 ;
		12'h839 : douta <= 12'h74D ;
		12'h83A : douta <= 12'h74A ;
		12'h83B : douta <= 12'h746 ;
		12'h83C : douta <= 12'h743 ;
		12'h83D : douta <= 12'h740 ;
		12'h83E : douta <= 12'h73D ;
		12'h83F : douta <= 12'h73A ;
		12'h840 : douta <= 12'h737 ;
		12'h841 : douta <= 12'h734 ;
		12'h842 : douta <= 12'h731 ;
		12'h843 : douta <= 12'h72D ;
		12'h844 : douta <= 12'h72A ;
		12'h845 : douta <= 12'h727 ;
		12'h846 : douta <= 12'h724 ;
		12'h847 : douta <= 12'h721 ;
		12'h848 : douta <= 12'h71E ;
		12'h849 : douta <= 12'h71B ;
		12'h84A : douta <= 12'h718 ;
		12'h84B : douta <= 12'h715 ;
		12'h84C : douta <= 12'h711 ;
		12'h84D : douta <= 12'h70E ;
		12'h84E : douta <= 12'h70B ;
		12'h84F : douta <= 12'h708 ;
		12'h850 : douta <= 12'h705 ;
		12'h851 : douta <= 12'h702 ;
		12'h852 : douta <= 12'h6FF ;
		12'h853 : douta <= 12'h6FC ;
		12'h854 : douta <= 12'h6F8 ;
		12'h855 : douta <= 12'h6F5 ;
		12'h856 : douta <= 12'h6F2 ;
		12'h857 : douta <= 12'h6EF ;
		12'h858 : douta <= 12'h6EC ;
		12'h859 : douta <= 12'h6E9 ;
		12'h85A : douta <= 12'h6E6 ;
		12'h85B : douta <= 12'h6E3 ;
		12'h85C : douta <= 12'h6E0 ;
		12'h85D : douta <= 12'h6DC ;
		12'h85E : douta <= 12'h6D9 ;
		12'h85F : douta <= 12'h6D6 ;
		12'h860 : douta <= 12'h6D3 ;
		12'h861 : douta <= 12'h6D0 ;
		12'h862 : douta <= 12'h6CD ;
		12'h863 : douta <= 12'h6CA ;
		12'h864 : douta <= 12'h6C7 ;
		12'h865 : douta <= 12'h6C4 ;
		12'h866 : douta <= 12'h6C1 ;
		12'h867 : douta <= 12'h6BD ;
		12'h868 : douta <= 12'h6BA ;
		12'h869 : douta <= 12'h6B7 ;
		12'h86A : douta <= 12'h6B4 ;
		12'h86B : douta <= 12'h6B1 ;
		12'h86C : douta <= 12'h6AE ;
		12'h86D : douta <= 12'h6AB ;
		12'h86E : douta <= 12'h6A8 ;
		12'h86F : douta <= 12'h6A5 ;
		12'h870 : douta <= 12'h6A2 ;
		12'h871 : douta <= 12'h69E ;
		12'h872 : douta <= 12'h69B ;
		12'h873 : douta <= 12'h698 ;
		12'h874 : douta <= 12'h695 ;
		12'h875 : douta <= 12'h692 ;
		12'h876 : douta <= 12'h68F ;
		12'h877 : douta <= 12'h68C ;
		12'h878 : douta <= 12'h689 ;
		12'h879 : douta <= 12'h686 ;
		12'h87A : douta <= 12'h683 ;
		12'h87B : douta <= 12'h680 ;
		12'h87C : douta <= 12'h67C ;
		12'h87D : douta <= 12'h679 ;
		12'h87E : douta <= 12'h676 ;
		12'h87F : douta <= 12'h673 ;
		12'h880 : douta <= 12'h670 ;
		12'h881 : douta <= 12'h66D ;
		12'h882 : douta <= 12'h66A ;
		12'h883 : douta <= 12'h667 ;
		12'h884 : douta <= 12'h664 ;
		12'h885 : douta <= 12'h661 ;
		12'h886 : douta <= 12'h65E ;
		12'h887 : douta <= 12'h65B ;
		12'h888 : douta <= 12'h658 ;
		12'h889 : douta <= 12'h654 ;
		12'h88A : douta <= 12'h651 ;
		12'h88B : douta <= 12'h64E ;
		12'h88C : douta <= 12'h64B ;
		12'h88D : douta <= 12'h648 ;
		12'h88E : douta <= 12'h645 ;
		12'h88F : douta <= 12'h642 ;
		12'h890 : douta <= 12'h63F ;
		12'h891 : douta <= 12'h63C ;
		12'h892 : douta <= 12'h639 ;
		12'h893 : douta <= 12'h636 ;
		12'h894 : douta <= 12'h633 ;
		12'h895 : douta <= 12'h630 ;
		12'h896 : douta <= 12'h62D ;
		12'h897 : douta <= 12'h62A ;
		12'h898 : douta <= 12'h627 ;
		12'h899 : douta <= 12'h623 ;
		12'h89A : douta <= 12'h620 ;
		12'h89B : douta <= 12'h61D ;
		12'h89C : douta <= 12'h61A ;
		12'h89D : douta <= 12'h617 ;
		12'h89E : douta <= 12'h614 ;
		12'h89F : douta <= 12'h611 ;
		12'h8A0 : douta <= 12'h60E ;
		12'h8A1 : douta <= 12'h60B ;
		12'h8A2 : douta <= 12'h608 ;
		12'h8A3 : douta <= 12'h605 ;
		12'h8A4 : douta <= 12'h602 ;
		12'h8A5 : douta <= 12'h5FF ;
		12'h8A6 : douta <= 12'h5FC ;
		12'h8A7 : douta <= 12'h5F9 ;
		12'h8A8 : douta <= 12'h5F6 ;
		12'h8A9 : douta <= 12'h5F3 ;
		12'h8AA : douta <= 12'h5F0 ;
		12'h8AB : douta <= 12'h5ED ;
		12'h8AC : douta <= 12'h5EA ;
		12'h8AD : douta <= 12'h5E7 ;
		12'h8AE : douta <= 12'h5E4 ;
		12'h8AF : douta <= 12'h5E1 ;
		12'h8B0 : douta <= 12'h5DE ;
		12'h8B1 : douta <= 12'h5DB ;
		12'h8B2 : douta <= 12'h5D7 ;
		12'h8B3 : douta <= 12'h5D4 ;
		12'h8B4 : douta <= 12'h5D1 ;
		12'h8B5 : douta <= 12'h5CE ;
		12'h8B6 : douta <= 12'h5CB ;
		12'h8B7 : douta <= 12'h5C8 ;
		12'h8B8 : douta <= 12'h5C5 ;
		12'h8B9 : douta <= 12'h5C2 ;
		12'h8BA : douta <= 12'h5BF ;
		12'h8BB : douta <= 12'h5BC ;
		12'h8BC : douta <= 12'h5B9 ;
		12'h8BD : douta <= 12'h5B6 ;
		12'h8BE : douta <= 12'h5B3 ;
		12'h8BF : douta <= 12'h5B0 ;
		12'h8C0 : douta <= 12'h5AD ;
		12'h8C1 : douta <= 12'h5AA ;
		12'h8C2 : douta <= 12'h5A7 ;
		12'h8C3 : douta <= 12'h5A4 ;
		12'h8C4 : douta <= 12'h5A1 ;
		12'h8C5 : douta <= 12'h59E ;
		12'h8C6 : douta <= 12'h59B ;
		12'h8C7 : douta <= 12'h598 ;
		12'h8C8 : douta <= 12'h595 ;
		12'h8C9 : douta <= 12'h592 ;
		12'h8CA : douta <= 12'h58F ;
		12'h8CB : douta <= 12'h58C ;
		12'h8CC : douta <= 12'h589 ;
		12'h8CD : douta <= 12'h586 ;
		12'h8CE : douta <= 12'h583 ;
		12'h8CF : douta <= 12'h580 ;
		12'h8D0 : douta <= 12'h57D ;
		12'h8D1 : douta <= 12'h57A ;
		12'h8D2 : douta <= 12'h577 ;
		12'h8D3 : douta <= 12'h574 ;
		12'h8D4 : douta <= 12'h571 ;
		12'h8D5 : douta <= 12'h56F ;
		12'h8D6 : douta <= 12'h56C ;
		12'h8D7 : douta <= 12'h569 ;
		12'h8D8 : douta <= 12'h566 ;
		12'h8D9 : douta <= 12'h563 ;
		12'h8DA : douta <= 12'h560 ;
		12'h8DB : douta <= 12'h55D ;
		12'h8DC : douta <= 12'h55A ;
		12'h8DD : douta <= 12'h557 ;
		12'h8DE : douta <= 12'h554 ;
		12'h8DF : douta <= 12'h551 ;
		12'h8E0 : douta <= 12'h54E ;
		12'h8E1 : douta <= 12'h54B ;
		12'h8E2 : douta <= 12'h548 ;
		12'h8E3 : douta <= 12'h545 ;
		12'h8E4 : douta <= 12'h542 ;
		12'h8E5 : douta <= 12'h53F ;
		12'h8E6 : douta <= 12'h53C ;
		12'h8E7 : douta <= 12'h539 ;
		12'h8E8 : douta <= 12'h536 ;
		12'h8E9 : douta <= 12'h533 ;
		12'h8EA : douta <= 12'h530 ;
		12'h8EB : douta <= 12'h52D ;
		12'h8EC : douta <= 12'h52B ;
		12'h8ED : douta <= 12'h528 ;
		12'h8EE : douta <= 12'h525 ;
		12'h8EF : douta <= 12'h522 ;
		12'h8F0 : douta <= 12'h51F ;
		12'h8F1 : douta <= 12'h51C ;
		12'h8F2 : douta <= 12'h519 ;
		12'h8F3 : douta <= 12'h516 ;
		12'h8F4 : douta <= 12'h513 ;
		12'h8F5 : douta <= 12'h510 ;
		12'h8F6 : douta <= 12'h50D ;
		12'h8F7 : douta <= 12'h50A ;
		12'h8F8 : douta <= 12'h507 ;
		12'h8F9 : douta <= 12'h504 ;
		12'h8FA : douta <= 12'h502 ;
		12'h8FB : douta <= 12'h4FF ;
		12'h8FC : douta <= 12'h4FC ;
		12'h8FD : douta <= 12'h4F9 ;
		12'h8FE : douta <= 12'h4F6 ;
		12'h8FF : douta <= 12'h4F3 ;
		12'h900 : douta <= 12'h4F0 ;
		12'h901 : douta <= 12'h4ED ;
		12'h902 : douta <= 12'h4EA ;
		12'h903 : douta <= 12'h4E7 ;
		12'h904 : douta <= 12'h4E5 ;
		12'h905 : douta <= 12'h4E2 ;
		12'h906 : douta <= 12'h4DF ;
		12'h907 : douta <= 12'h4DC ;
		12'h908 : douta <= 12'h4D9 ;
		12'h909 : douta <= 12'h4D6 ;
		12'h90A : douta <= 12'h4D3 ;
		12'h90B : douta <= 12'h4D0 ;
		12'h90C : douta <= 12'h4CD ;
		12'h90D : douta <= 12'h4CB ;
		12'h90E : douta <= 12'h4C8 ;
		12'h90F : douta <= 12'h4C5 ;
		12'h910 : douta <= 12'h4C2 ;
		12'h911 : douta <= 12'h4BF ;
		12'h912 : douta <= 12'h4BC ;
		12'h913 : douta <= 12'h4B9 ;
		12'h914 : douta <= 12'h4B7 ;
		12'h915 : douta <= 12'h4B4 ;
		12'h916 : douta <= 12'h4B1 ;
		12'h917 : douta <= 12'h4AE ;
		12'h918 : douta <= 12'h4AB ;
		12'h919 : douta <= 12'h4A8 ;
		12'h91A : douta <= 12'h4A5 ;
		12'h91B : douta <= 12'h4A3 ;
		12'h91C : douta <= 12'h4A0 ;
		12'h91D : douta <= 12'h49D ;
		12'h91E : douta <= 12'h49A ;
		12'h91F : douta <= 12'h497 ;
		12'h920 : douta <= 12'h494 ;
		12'h921 : douta <= 12'h491 ;
		12'h922 : douta <= 12'h48F ;
		12'h923 : douta <= 12'h48C ;
		12'h924 : douta <= 12'h489 ;
		12'h925 : douta <= 12'h486 ;
		12'h926 : douta <= 12'h483 ;
		12'h927 : douta <= 12'h480 ;
		12'h928 : douta <= 12'h47E ;
		12'h929 : douta <= 12'h47B ;
		12'h92A : douta <= 12'h478 ;
		12'h92B : douta <= 12'h475 ;
		12'h92C : douta <= 12'h472 ;
		12'h92D : douta <= 12'h470 ;
		12'h92E : douta <= 12'h46D ;
		12'h92F : douta <= 12'h46A ;
		12'h930 : douta <= 12'h467 ;
		12'h931 : douta <= 12'h464 ;
		12'h932 : douta <= 12'h462 ;
		12'h933 : douta <= 12'h45F ;
		12'h934 : douta <= 12'h45C ;
		12'h935 : douta <= 12'h459 ;
		12'h936 : douta <= 12'h456 ;
		12'h937 : douta <= 12'h454 ;
		12'h938 : douta <= 12'h451 ;
		12'h939 : douta <= 12'h44E ;
		12'h93A : douta <= 12'h44B ;
		12'h93B : douta <= 12'h448 ;
		12'h93C : douta <= 12'h446 ;
		12'h93D : douta <= 12'h443 ;
		12'h93E : douta <= 12'h440 ;
		12'h93F : douta <= 12'h43D ;
		12'h940 : douta <= 12'h43B ;
		12'h941 : douta <= 12'h438 ;
		12'h942 : douta <= 12'h435 ;
		12'h943 : douta <= 12'h432 ;
		12'h944 : douta <= 12'h42F ;
		12'h945 : douta <= 12'h42D ;
		12'h946 : douta <= 12'h42A ;
		12'h947 : douta <= 12'h427 ;
		12'h948 : douta <= 12'h424 ;
		12'h949 : douta <= 12'h422 ;
		12'h94A : douta <= 12'h41F ;
		12'h94B : douta <= 12'h41C ;
		12'h94C : douta <= 12'h419 ;
		12'h94D : douta <= 12'h417 ;
		12'h94E : douta <= 12'h414 ;
		12'h94F : douta <= 12'h411 ;
		12'h950 : douta <= 12'h40F ;
		12'h951 : douta <= 12'h40C ;
		12'h952 : douta <= 12'h409 ;
		12'h953 : douta <= 12'h406 ;
		12'h954 : douta <= 12'h404 ;
		12'h955 : douta <= 12'h401 ;
		12'h956 : douta <= 12'h3FE ;
		12'h957 : douta <= 12'h3FB ;
		12'h958 : douta <= 12'h3F9 ;
		12'h959 : douta <= 12'h3F6 ;
		12'h95A : douta <= 12'h3F3 ;
		12'h95B : douta <= 12'h3F1 ;
		12'h95C : douta <= 12'h3EE ;
		12'h95D : douta <= 12'h3EB ;
		12'h95E : douta <= 12'h3E9 ;
		12'h95F : douta <= 12'h3E6 ;
		12'h960 : douta <= 12'h3E3 ;
		12'h961 : douta <= 12'h3E0 ;
		12'h962 : douta <= 12'h3DE ;
		12'h963 : douta <= 12'h3DB ;
		12'h964 : douta <= 12'h3D8 ;
		12'h965 : douta <= 12'h3D6 ;
		12'h966 : douta <= 12'h3D3 ;
		12'h967 : douta <= 12'h3D0 ;
		12'h968 : douta <= 12'h3CE ;
		12'h969 : douta <= 12'h3CB ;
		12'h96A : douta <= 12'h3C8 ;
		12'h96B : douta <= 12'h3C6 ;
		12'h96C : douta <= 12'h3C3 ;
		12'h96D : douta <= 12'h3C0 ;
		12'h96E : douta <= 12'h3BE ;
		12'h96F : douta <= 12'h3BB ;
		12'h970 : douta <= 12'h3B8 ;
		12'h971 : douta <= 12'h3B6 ;
		12'h972 : douta <= 12'h3B3 ;
		12'h973 : douta <= 12'h3B0 ;
		12'h974 : douta <= 12'h3AE ;
		12'h975 : douta <= 12'h3AB ;
		12'h976 : douta <= 12'h3A8 ;
		12'h977 : douta <= 12'h3A6 ;
		12'h978 : douta <= 12'h3A3 ;
		12'h979 : douta <= 12'h3A1 ;
		12'h97A : douta <= 12'h39E ;
		12'h97B : douta <= 12'h39B ;
		12'h97C : douta <= 12'h399 ;
		12'h97D : douta <= 12'h396 ;
		12'h97E : douta <= 12'h393 ;
		12'h97F : douta <= 12'h391 ;
		12'h980 : douta <= 12'h38E ;
		12'h981 : douta <= 12'h38C ;
		12'h982 : douta <= 12'h389 ;
		12'h983 : douta <= 12'h386 ;
		12'h984 : douta <= 12'h384 ;
		12'h985 : douta <= 12'h381 ;
		12'h986 : douta <= 12'h37F ;
		12'h987 : douta <= 12'h37C ;
		12'h988 : douta <= 12'h379 ;
		12'h989 : douta <= 12'h377 ;
		12'h98A : douta <= 12'h374 ;
		12'h98B : douta <= 12'h372 ;
		12'h98C : douta <= 12'h36F ;
		12'h98D : douta <= 12'h36D ;
		12'h98E : douta <= 12'h36A ;
		12'h98F : douta <= 12'h367 ;
		12'h990 : douta <= 12'h365 ;
		12'h991 : douta <= 12'h362 ;
		12'h992 : douta <= 12'h360 ;
		12'h993 : douta <= 12'h35D ;
		12'h994 : douta <= 12'h35B ;
		12'h995 : douta <= 12'h358 ;
		12'h996 : douta <= 12'h355 ;
		12'h997 : douta <= 12'h353 ;
		12'h998 : douta <= 12'h350 ;
		12'h999 : douta <= 12'h34E ;
		12'h99A : douta <= 12'h34B ;
		12'h99B : douta <= 12'h349 ;
		12'h99C : douta <= 12'h346 ;
		12'h99D : douta <= 12'h344 ;
		12'h99E : douta <= 12'h341 ;
		12'h99F : douta <= 12'h33F ;
		12'h9A0 : douta <= 12'h33C ;
		12'h9A1 : douta <= 12'h33A ;
		12'h9A2 : douta <= 12'h337 ;
		12'h9A3 : douta <= 12'h335 ;
		12'h9A4 : douta <= 12'h332 ;
		12'h9A5 : douta <= 12'h330 ;
		12'h9A6 : douta <= 12'h32D ;
		12'h9A7 : douta <= 12'h32B ;
		12'h9A8 : douta <= 12'h328 ;
		12'h9A9 : douta <= 12'h326 ;
		12'h9AA : douta <= 12'h323 ;
		12'h9AB : douta <= 12'h321 ;
		12'h9AC : douta <= 12'h31E ;
		12'h9AD : douta <= 12'h31C ;
		12'h9AE : douta <= 12'h319 ;
		12'h9AF : douta <= 12'h317 ;
		12'h9B0 : douta <= 12'h314 ;
		12'h9B1 : douta <= 12'h312 ;
		12'h9B2 : douta <= 12'h30F ;
		12'h9B3 : douta <= 12'h30D ;
		12'h9B4 : douta <= 12'h30A ;
		12'h9B5 : douta <= 12'h308 ;
		12'h9B6 : douta <= 12'h305 ;
		12'h9B7 : douta <= 12'h303 ;
		12'h9B8 : douta <= 12'h300 ;
		12'h9B9 : douta <= 12'h2FE ;
		12'h9BA : douta <= 12'h2FC ;
		12'h9BB : douta <= 12'h2F9 ;
		12'h9BC : douta <= 12'h2F7 ;
		12'h9BD : douta <= 12'h2F4 ;
		12'h9BE : douta <= 12'h2F2 ;
		12'h9BF : douta <= 12'h2EF ;
		12'h9C0 : douta <= 12'h2ED ;
		12'h9C1 : douta <= 12'h2EA ;
		12'h9C2 : douta <= 12'h2E8 ;
		12'h9C3 : douta <= 12'h2E6 ;
		12'h9C4 : douta <= 12'h2E3 ;
		12'h9C5 : douta <= 12'h2E1 ;
		12'h9C6 : douta <= 12'h2DE ;
		12'h9C7 : douta <= 12'h2DC ;
		12'h9C8 : douta <= 12'h2DA ;
		12'h9C9 : douta <= 12'h2D7 ;
		12'h9CA : douta <= 12'h2D5 ;
		12'h9CB : douta <= 12'h2D2 ;
		12'h9CC : douta <= 12'h2D0 ;
		12'h9CD : douta <= 12'h2CE ;
		12'h9CE : douta <= 12'h2CB ;
		12'h9CF : douta <= 12'h2C9 ;
		12'h9D0 : douta <= 12'h2C6 ;
		12'h9D1 : douta <= 12'h2C4 ;
		12'h9D2 : douta <= 12'h2C2 ;
		12'h9D3 : douta <= 12'h2BF ;
		12'h9D4 : douta <= 12'h2BD ;
		12'h9D5 : douta <= 12'h2BB ;
		12'h9D6 : douta <= 12'h2B8 ;
		12'h9D7 : douta <= 12'h2B6 ;
		12'h9D8 : douta <= 12'h2B4 ;
		12'h9D9 : douta <= 12'h2B1 ;
		12'h9DA : douta <= 12'h2AF ;
		12'h9DB : douta <= 12'h2AC ;
		12'h9DC : douta <= 12'h2AA ;
		12'h9DD : douta <= 12'h2A8 ;
		12'h9DE : douta <= 12'h2A5 ;
		12'h9DF : douta <= 12'h2A3 ;
		12'h9E0 : douta <= 12'h2A1 ;
		12'h9E1 : douta <= 12'h29E ;
		12'h9E2 : douta <= 12'h29C ;
		12'h9E3 : douta <= 12'h29A ;
		12'h9E4 : douta <= 12'h298 ;
		12'h9E5 : douta <= 12'h295 ;
		12'h9E6 : douta <= 12'h293 ;
		12'h9E7 : douta <= 12'h291 ;
		12'h9E8 : douta <= 12'h28E ;
		12'h9E9 : douta <= 12'h28C ;
		12'h9EA : douta <= 12'h28A ;
		12'h9EB : douta <= 12'h287 ;
		12'h9EC : douta <= 12'h285 ;
		12'h9ED : douta <= 12'h283 ;
		12'h9EE : douta <= 12'h281 ;
		12'h9EF : douta <= 12'h27E ;
		12'h9F0 : douta <= 12'h27C ;
		12'h9F1 : douta <= 12'h27A ;
		12'h9F2 : douta <= 12'h277 ;
		12'h9F3 : douta <= 12'h275 ;
		12'h9F4 : douta <= 12'h273 ;
		12'h9F5 : douta <= 12'h271 ;
		12'h9F6 : douta <= 12'h26E ;
		12'h9F7 : douta <= 12'h26C ;
		12'h9F8 : douta <= 12'h26A ;
		12'h9F9 : douta <= 12'h268 ;
		12'h9FA : douta <= 12'h265 ;
		12'h9FB : douta <= 12'h263 ;
		12'h9FC : douta <= 12'h261 ;
		12'h9FD : douta <= 12'h25F ;
		12'h9FE : douta <= 12'h25C ;
		12'h9FF : douta <= 12'h25A ;
		12'hA00 : douta <= 12'h258 ;
		12'hA01 : douta <= 12'h256 ;
		12'hA02 : douta <= 12'h254 ;
		12'hA03 : douta <= 12'h251 ;
		12'hA04 : douta <= 12'h24F ;
		12'hA05 : douta <= 12'h24D ;
		12'hA06 : douta <= 12'h24B ;
		12'hA07 : douta <= 12'h249 ;
		12'hA08 : douta <= 12'h246 ;
		12'hA09 : douta <= 12'h244 ;
		12'hA0A : douta <= 12'h242 ;
		12'hA0B : douta <= 12'h240 ;
		12'hA0C : douta <= 12'h23E ;
		12'hA0D : douta <= 12'h23B ;
		12'hA0E : douta <= 12'h239 ;
		12'hA0F : douta <= 12'h237 ;
		12'hA10 : douta <= 12'h235 ;
		12'hA11 : douta <= 12'h233 ;
		12'hA12 : douta <= 12'h231 ;
		12'hA13 : douta <= 12'h22E ;
		12'hA14 : douta <= 12'h22C ;
		12'hA15 : douta <= 12'h22A ;
		12'hA16 : douta <= 12'h228 ;
		12'hA17 : douta <= 12'h226 ;
		12'hA18 : douta <= 12'h224 ;
		12'hA19 : douta <= 12'h222 ;
		12'hA1A : douta <= 12'h21F ;
		12'hA1B : douta <= 12'h21D ;
		12'hA1C : douta <= 12'h21B ;
		12'hA1D : douta <= 12'h219 ;
		12'hA1E : douta <= 12'h217 ;
		12'hA1F : douta <= 12'h215 ;
		12'hA20 : douta <= 12'h213 ;
		12'hA21 : douta <= 12'h211 ;
		12'hA22 : douta <= 12'h20F ;
		12'hA23 : douta <= 12'h20C ;
		12'hA24 : douta <= 12'h20A ;
		12'hA25 : douta <= 12'h208 ;
		12'hA26 : douta <= 12'h206 ;
		12'hA27 : douta <= 12'h204 ;
		12'hA28 : douta <= 12'h202 ;
		12'hA29 : douta <= 12'h200 ;
		12'hA2A : douta <= 12'h1FE ;
		12'hA2B : douta <= 12'h1FC ;
		12'hA2C : douta <= 12'h1FA ;
		12'hA2D : douta <= 12'h1F8 ;
		12'hA2E : douta <= 12'h1F6 ;
		12'hA2F : douta <= 12'h1F4 ;
		12'hA30 : douta <= 12'h1F1 ;
		12'hA31 : douta <= 12'h1EF ;
		12'hA32 : douta <= 12'h1ED ;
		12'hA33 : douta <= 12'h1EB ;
		12'hA34 : douta <= 12'h1E9 ;
		12'hA35 : douta <= 12'h1E7 ;
		12'hA36 : douta <= 12'h1E5 ;
		12'hA37 : douta <= 12'h1E3 ;
		12'hA38 : douta <= 12'h1E1 ;
		12'hA39 : douta <= 12'h1DF ;
		12'hA3A : douta <= 12'h1DD ;
		12'hA3B : douta <= 12'h1DB ;
		12'hA3C : douta <= 12'h1D9 ;
		12'hA3D : douta <= 12'h1D7 ;
		12'hA3E : douta <= 12'h1D5 ;
		12'hA3F : douta <= 12'h1D3 ;
		12'hA40 : douta <= 12'h1D1 ;
		12'hA41 : douta <= 12'h1CF ;
		12'hA42 : douta <= 12'h1CD ;
		12'hA43 : douta <= 12'h1CB ;
		12'hA44 : douta <= 12'h1C9 ;
		12'hA45 : douta <= 12'h1C7 ;
		12'hA46 : douta <= 12'h1C5 ;
		12'hA47 : douta <= 12'h1C3 ;
		12'hA48 : douta <= 12'h1C1 ;
		12'hA49 : douta <= 12'h1BF ;
		12'hA4A : douta <= 12'h1BD ;
		12'hA4B : douta <= 12'h1BB ;
		12'hA4C : douta <= 12'h1BA ;
		12'hA4D : douta <= 12'h1B8 ;
		12'hA4E : douta <= 12'h1B6 ;
		12'hA4F : douta <= 12'h1B4 ;
		12'hA50 : douta <= 12'h1B2 ;
		12'hA51 : douta <= 12'h1B0 ;
		12'hA52 : douta <= 12'h1AE ;
		12'hA53 : douta <= 12'h1AC ;
		12'hA54 : douta <= 12'h1AA ;
		12'hA55 : douta <= 12'h1A8 ;
		12'hA56 : douta <= 12'h1A6 ;
		12'hA57 : douta <= 12'h1A4 ;
		12'hA58 : douta <= 12'h1A2 ;
		12'hA59 : douta <= 12'h1A1 ;
		12'hA5A : douta <= 12'h19F ;
		12'hA5B : douta <= 12'h19D ;
		12'hA5C : douta <= 12'h19B ;
		12'hA5D : douta <= 12'h199 ;
		12'hA5E : douta <= 12'h197 ;
		12'hA5F : douta <= 12'h195 ;
		12'hA60 : douta <= 12'h193 ;
		12'hA61 : douta <= 12'h191 ;
		12'hA62 : douta <= 12'h190 ;
		12'hA63 : douta <= 12'h18E ;
		12'hA64 : douta <= 12'h18C ;
		12'hA65 : douta <= 12'h18A ;
		12'hA66 : douta <= 12'h188 ;
		12'hA67 : douta <= 12'h186 ;
		12'hA68 : douta <= 12'h184 ;
		12'hA69 : douta <= 12'h183 ;
		12'hA6A : douta <= 12'h181 ;
		12'hA6B : douta <= 12'h17F ;
		12'hA6C : douta <= 12'h17D ;
		12'hA6D : douta <= 12'h17B ;
		12'hA6E : douta <= 12'h17A ;
		12'hA6F : douta <= 12'h178 ;
		12'hA70 : douta <= 12'h176 ;
		12'hA71 : douta <= 12'h174 ;
		12'hA72 : douta <= 12'h172 ;
		12'hA73 : douta <= 12'h170 ;
		12'hA74 : douta <= 12'h16F ;
		12'hA75 : douta <= 12'h16D ;
		12'hA76 : douta <= 12'h16B ;
		12'hA77 : douta <= 12'h169 ;
		12'hA78 : douta <= 12'h168 ;
		12'hA79 : douta <= 12'h166 ;
		12'hA7A : douta <= 12'h164 ;
		12'hA7B : douta <= 12'h162 ;
		12'hA7C : douta <= 12'h160 ;
		12'hA7D : douta <= 12'h15F ;
		12'hA7E : douta <= 12'h15D ;
		12'hA7F : douta <= 12'h15B ;
		12'hA80 : douta <= 12'h159 ;
		12'hA81 : douta <= 12'h158 ;
		12'hA82 : douta <= 12'h156 ;
		12'hA83 : douta <= 12'h154 ;
		12'hA84 : douta <= 12'h153 ;
		12'hA85 : douta <= 12'h151 ;
		12'hA86 : douta <= 12'h14F ;
		12'hA87 : douta <= 12'h14D ;
		12'hA88 : douta <= 12'h14C ;
		12'hA89 : douta <= 12'h14A ;
		12'hA8A : douta <= 12'h148 ;
		12'hA8B : douta <= 12'h147 ;
		12'hA8C : douta <= 12'h145 ;
		12'hA8D : douta <= 12'h143 ;
		12'hA8E : douta <= 12'h141 ;
		12'hA8F : douta <= 12'h140 ;
		12'hA90 : douta <= 12'h13E ;
		12'hA91 : douta <= 12'h13C ;
		12'hA92 : douta <= 12'h13B ;
		12'hA93 : douta <= 12'h139 ;
		12'hA94 : douta <= 12'h137 ;
		12'hA95 : douta <= 12'h136 ;
		12'hA96 : douta <= 12'h134 ;
		12'hA97 : douta <= 12'h132 ;
		12'hA98 : douta <= 12'h131 ;
		12'hA99 : douta <= 12'h12F ;
		12'hA9A : douta <= 12'h12D ;
		12'hA9B : douta <= 12'h12C ;
		12'hA9C : douta <= 12'h12A ;
		12'hA9D : douta <= 12'h129 ;
		12'hA9E : douta <= 12'h127 ;
		12'hA9F : douta <= 12'h125 ;
		12'hAA0 : douta <= 12'h124 ;
		12'hAA1 : douta <= 12'h122 ;
		12'hAA2 : douta <= 12'h121 ;
		12'hAA3 : douta <= 12'h11F ;
		12'hAA4 : douta <= 12'h11D ;
		12'hAA5 : douta <= 12'h11C ;
		12'hAA6 : douta <= 12'h11A ;
		12'hAA7 : douta <= 12'h119 ;
		12'hAA8 : douta <= 12'h117 ;
		12'hAA9 : douta <= 12'h115 ;
		12'hAAA : douta <= 12'h114 ;
		12'hAAB : douta <= 12'h112 ;
		12'hAAC : douta <= 12'h111 ;
		12'hAAD : douta <= 12'h10F ;
		12'hAAE : douta <= 12'h10E ;
		12'hAAF : douta <= 12'h10C ;
		12'hAB0 : douta <= 12'h10A ;
		12'hAB1 : douta <= 12'h109 ;
		12'hAB2 : douta <= 12'h107 ;
		12'hAB3 : douta <= 12'h106 ;
		12'hAB4 : douta <= 12'h104 ;
		12'hAB5 : douta <= 12'h103 ;
		12'hAB6 : douta <= 12'h101 ;
		12'hAB7 : douta <= 12'h100 ;
		12'hAB8 : douta <= 12'h0FE ;
		12'hAB9 : douta <= 12'h0FD ;
		12'hABA : douta <= 12'h0FB ;
		12'hABB : douta <= 12'h0FA ;
		12'hABC : douta <= 12'h0F8 ;
		12'hABD : douta <= 12'h0F7 ;
		12'hABE : douta <= 12'h0F5 ;
		12'hABF : douta <= 12'h0F4 ;
		12'hAC0 : douta <= 12'h0F2 ;
		12'hAC1 : douta <= 12'h0F1 ;
		12'hAC2 : douta <= 12'h0EF ;
		12'hAC3 : douta <= 12'h0EE ;
		12'hAC4 : douta <= 12'h0EC ;
		12'hAC5 : douta <= 12'h0EB ;
		12'hAC6 : douta <= 12'h0E9 ;
		12'hAC7 : douta <= 12'h0E8 ;
		12'hAC8 : douta <= 12'h0E7 ;
		12'hAC9 : douta <= 12'h0E5 ;
		12'hACA : douta <= 12'h0E4 ;
		12'hACB : douta <= 12'h0E2 ;
		12'hACC : douta <= 12'h0E1 ;
		12'hACD : douta <= 12'h0DF ;
		12'hACE : douta <= 12'h0DE ;
		12'hACF : douta <= 12'h0DC ;
		12'hAD0 : douta <= 12'h0DB ;
		12'hAD1 : douta <= 12'h0DA ;
		12'hAD2 : douta <= 12'h0D8 ;
		12'hAD3 : douta <= 12'h0D7 ;
		12'hAD4 : douta <= 12'h0D5 ;
		12'hAD5 : douta <= 12'h0D4 ;
		12'hAD6 : douta <= 12'h0D3 ;
		12'hAD7 : douta <= 12'h0D1 ;
		12'hAD8 : douta <= 12'h0D0 ;
		12'hAD9 : douta <= 12'h0CF ;
		12'hADA : douta <= 12'h0CD ;
		12'hADB : douta <= 12'h0CC ;
		12'hADC : douta <= 12'h0CA ;
		12'hADD : douta <= 12'h0C9 ;
		12'hADE : douta <= 12'h0C8 ;
		12'hADF : douta <= 12'h0C6 ;
		12'hAE0 : douta <= 12'h0C5 ;
		12'hAE1 : douta <= 12'h0C4 ;
		12'hAE2 : douta <= 12'h0C2 ;
		12'hAE3 : douta <= 12'h0C1 ;
		12'hAE4 : douta <= 12'h0C0 ;
		12'hAE5 : douta <= 12'h0BE ;
		12'hAE6 : douta <= 12'h0BD ;
		12'hAE7 : douta <= 12'h0BC ;
		12'hAE8 : douta <= 12'h0BA ;
		12'hAE9 : douta <= 12'h0B9 ;
		12'hAEA : douta <= 12'h0B8 ;
		12'hAEB : douta <= 12'h0B7 ;
		12'hAEC : douta <= 12'h0B5 ;
		12'hAED : douta <= 12'h0B4 ;
		12'hAEE : douta <= 12'h0B3 ;
		12'hAEF : douta <= 12'h0B1 ;
		12'hAF0 : douta <= 12'h0B0 ;
		12'hAF1 : douta <= 12'h0AF ;
		12'hAF2 : douta <= 12'h0AE ;
		12'hAF3 : douta <= 12'h0AC ;
		12'hAF4 : douta <= 12'h0AB ;
		12'hAF5 : douta <= 12'h0AA ;
		12'hAF6 : douta <= 12'h0A9 ;
		12'hAF7 : douta <= 12'h0A7 ;
		12'hAF8 : douta <= 12'h0A6 ;
		12'hAF9 : douta <= 12'h0A5 ;
		12'hAFA : douta <= 12'h0A4 ;
		12'hAFB : douta <= 12'h0A2 ;
		12'hAFC : douta <= 12'h0A1 ;
		12'hAFD : douta <= 12'h0A0 ;
		12'hAFE : douta <= 12'h09F ;
		12'hAFF : douta <= 12'h09E ;
		12'hB00 : douta <= 12'h09C ;
		12'hB01 : douta <= 12'h09B ;
		12'hB02 : douta <= 12'h09A ;
		12'hB03 : douta <= 12'h099 ;
		12'hB04 : douta <= 12'h098 ;
		12'hB05 : douta <= 12'h096 ;
		12'hB06 : douta <= 12'h095 ;
		12'hB07 : douta <= 12'h094 ;
		12'hB08 : douta <= 12'h093 ;
		12'hB09 : douta <= 12'h092 ;
		12'hB0A : douta <= 12'h091 ;
		12'hB0B : douta <= 12'h08F ;
		12'hB0C : douta <= 12'h08E ;
		12'hB0D : douta <= 12'h08D ;
		12'hB0E : douta <= 12'h08C ;
		12'hB0F : douta <= 12'h08B ;
		12'hB10 : douta <= 12'h08A ;
		12'hB11 : douta <= 12'h089 ;
		12'hB12 : douta <= 12'h087 ;
		12'hB13 : douta <= 12'h086 ;
		12'hB14 : douta <= 12'h085 ;
		12'hB15 : douta <= 12'h084 ;
		12'hB16 : douta <= 12'h083 ;
		12'hB17 : douta <= 12'h082 ;
		12'hB18 : douta <= 12'h081 ;
		12'hB19 : douta <= 12'h080 ;
		12'hB1A : douta <= 12'h07F ;
		12'hB1B : douta <= 12'h07E ;
		12'hB1C : douta <= 12'h07C ;
		12'hB1D : douta <= 12'h07B ;
		12'hB1E : douta <= 12'h07A ;
		12'hB1F : douta <= 12'h079 ;
		12'hB20 : douta <= 12'h078 ;
		12'hB21 : douta <= 12'h077 ;
		12'hB22 : douta <= 12'h076 ;
		12'hB23 : douta <= 12'h075 ;
		12'hB24 : douta <= 12'h074 ;
		12'hB25 : douta <= 12'h073 ;
		12'hB26 : douta <= 12'h072 ;
		12'hB27 : douta <= 12'h071 ;
		12'hB28 : douta <= 12'h070 ;
		12'hB29 : douta <= 12'h06F ;
		12'hB2A : douta <= 12'h06E ;
		12'hB2B : douta <= 12'h06D ;
		12'hB2C : douta <= 12'h06C ;
		12'hB2D : douta <= 12'h06B ;
		12'hB2E : douta <= 12'h06A ;
		12'hB2F : douta <= 12'h069 ;
		12'hB30 : douta <= 12'h068 ;
		12'hB31 : douta <= 12'h067 ;
		12'hB32 : douta <= 12'h066 ;
		12'hB33 : douta <= 12'h065 ;
		12'hB34 : douta <= 12'h064 ;
		12'hB35 : douta <= 12'h063 ;
		12'hB36 : douta <= 12'h062 ;
		12'hB37 : douta <= 12'h061 ;
		12'hB38 : douta <= 12'h060 ;
		12'hB39 : douta <= 12'h05F ;
		12'hB3A : douta <= 12'h05E ;
		12'hB3B : douta <= 12'h05D ;
		12'hB3C : douta <= 12'h05C ;
		12'hB3D : douta <= 12'h05B ;
		12'hB3E : douta <= 12'h05A ;
		12'hB3F : douta <= 12'h05A ;
		12'hB40 : douta <= 12'h059 ;
		12'hB41 : douta <= 12'h058 ;
		12'hB42 : douta <= 12'h057 ;
		12'hB43 : douta <= 12'h056 ;
		12'hB44 : douta <= 12'h055 ;
		12'hB45 : douta <= 12'h054 ;
		12'hB46 : douta <= 12'h053 ;
		12'hB47 : douta <= 12'h052 ;
		12'hB48 : douta <= 12'h051 ;
		12'hB49 : douta <= 12'h051 ;
		12'hB4A : douta <= 12'h050 ;
		12'hB4B : douta <= 12'h04F ;
		12'hB4C : douta <= 12'h04E ;
		12'hB4D : douta <= 12'h04D ;
		12'hB4E : douta <= 12'h04C ;
		12'hB4F : douta <= 12'h04B ;
		12'hB50 : douta <= 12'h04B ;
		12'hB51 : douta <= 12'h04A ;
		12'hB52 : douta <= 12'h049 ;
		12'hB53 : douta <= 12'h048 ;
		12'hB54 : douta <= 12'h047 ;
		12'hB55 : douta <= 12'h047 ;
		12'hB56 : douta <= 12'h046 ;
		12'hB57 : douta <= 12'h045 ;
		12'hB58 : douta <= 12'h044 ;
		12'hB59 : douta <= 12'h043 ;
		12'hB5A : douta <= 12'h043 ;
		12'hB5B : douta <= 12'h042 ;
		12'hB5C : douta <= 12'h041 ;
		12'hB5D : douta <= 12'h040 ;
		12'hB5E : douta <= 12'h03F ;
		12'hB5F : douta <= 12'h03F ;
		12'hB60 : douta <= 12'h03E ;
		12'hB61 : douta <= 12'h03D ;
		12'hB62 : douta <= 12'h03C ;
		12'hB63 : douta <= 12'h03C ;
		12'hB64 : douta <= 12'h03B ;
		12'hB65 : douta <= 12'h03A ;
		12'hB66 : douta <= 12'h039 ;
		12'hB67 : douta <= 12'h039 ;
		12'hB68 : douta <= 12'h038 ;
		12'hB69 : douta <= 12'h037 ;
		12'hB6A : douta <= 12'h036 ;
		12'hB6B : douta <= 12'h036 ;
		12'hB6C : douta <= 12'h035 ;
		12'hB6D : douta <= 12'h034 ;
		12'hB6E : douta <= 12'h034 ;
		12'hB6F : douta <= 12'h033 ;
		12'hB70 : douta <= 12'h032 ;
		12'hB71 : douta <= 12'h032 ;
		12'hB72 : douta <= 12'h031 ;
		12'hB73 : douta <= 12'h030 ;
		12'hB74 : douta <= 12'h030 ;
		12'hB75 : douta <= 12'h02F ;
		12'hB76 : douta <= 12'h02E ;
		12'hB77 : douta <= 12'h02E ;
		12'hB78 : douta <= 12'h02D ;
		12'hB79 : douta <= 12'h02C ;
		12'hB7A : douta <= 12'h02C ;
		12'hB7B : douta <= 12'h02B ;
		12'hB7C : douta <= 12'h02A ;
		12'hB7D : douta <= 12'h02A ;
		12'hB7E : douta <= 12'h029 ;
		12'hB7F : douta <= 12'h028 ;
		12'hB80 : douta <= 12'h028 ;
		12'hB81 : douta <= 12'h027 ;
		12'hB82 : douta <= 12'h027 ;
		12'hB83 : douta <= 12'h026 ;
		12'hB84 : douta <= 12'h025 ;
		12'hB85 : douta <= 12'h025 ;
		12'hB86 : douta <= 12'h024 ;
		12'hB87 : douta <= 12'h024 ;
		12'hB88 : douta <= 12'h023 ;
		12'hB89 : douta <= 12'h023 ;
		12'hB8A : douta <= 12'h022 ;
		12'hB8B : douta <= 12'h021 ;
		12'hB8C : douta <= 12'h021 ;
		12'hB8D : douta <= 12'h020 ;
		12'hB8E : douta <= 12'h020 ;
		12'hB8F : douta <= 12'h01F ;
		12'hB90 : douta <= 12'h01F ;
		12'hB91 : douta <= 12'h01E ;
		12'hB92 : douta <= 12'h01E ;
		12'hB93 : douta <= 12'h01D ;
		12'hB94 : douta <= 12'h01D ;
		12'hB95 : douta <= 12'h01C ;
		12'hB96 : douta <= 12'h01C ;
		12'hB97 : douta <= 12'h01B ;
		12'hB98 : douta <= 12'h01A ;
		12'hB99 : douta <= 12'h01A ;
		12'hB9A : douta <= 12'h01A ;
		12'hB9B : douta <= 12'h019 ;
		12'hB9C : douta <= 12'h019 ;
		12'hB9D : douta <= 12'h018 ;
		12'hB9E : douta <= 12'h018 ;
		12'hB9F : douta <= 12'h017 ;
		12'hBA0 : douta <= 12'h017 ;
		12'hBA1 : douta <= 12'h016 ;
		12'hBA2 : douta <= 12'h016 ;
		12'hBA3 : douta <= 12'h015 ;
		12'hBA4 : douta <= 12'h015 ;
		12'hBA5 : douta <= 12'h014 ;
		12'hBA6 : douta <= 12'h014 ;
		12'hBA7 : douta <= 12'h014 ;
		12'hBA8 : douta <= 12'h013 ;
		12'hBA9 : douta <= 12'h013 ;
		12'hBAA : douta <= 12'h012 ;
		12'hBAB : douta <= 12'h012 ;
		12'hBAC : douta <= 12'h011 ;
		12'hBAD : douta <= 12'h011 ;
		12'hBAE : douta <= 12'h011 ;
		12'hBAF : douta <= 12'h010 ;
		12'hBB0 : douta <= 12'h010 ;
		12'hBB1 : douta <= 12'h010 ;
		12'hBB2 : douta <= 12'h00F ;
		12'hBB3 : douta <= 12'h00F ;
		12'hBB4 : douta <= 12'h00E ;
		12'hBB5 : douta <= 12'h00E ;
		12'hBB6 : douta <= 12'h00E ;
		12'hBB7 : douta <= 12'h00D ;
		12'hBB8 : douta <= 12'h00D ;
		12'hBB9 : douta <= 12'h00D ;
		12'hBBA : douta <= 12'h00C ;
		12'hBBB : douta <= 12'h00C ;
		12'hBBC : douta <= 12'h00C ;
		12'hBBD : douta <= 12'h00B ;
		12'hBBE : douta <= 12'h00B ;
		12'hBBF : douta <= 12'h00B ;
		12'hBC0 : douta <= 12'h00A ;
		12'hBC1 : douta <= 12'h00A ;
		12'hBC2 : douta <= 12'h00A ;
		12'hBC3 : douta <= 12'h009 ;
		12'hBC4 : douta <= 12'h009 ;
		12'hBC5 : douta <= 12'h009 ;
		12'hBC6 : douta <= 12'h009 ;
		12'hBC7 : douta <= 12'h008 ;
		12'hBC8 : douta <= 12'h008 ;
		12'hBC9 : douta <= 12'h008 ;
		12'hBCA : douta <= 12'h008 ;
		12'hBCB : douta <= 12'h007 ;
		12'hBCC : douta <= 12'h007 ;
		12'hBCD : douta <= 12'h007 ;
		12'hBCE : douta <= 12'h007 ;
		12'hBCF : douta <= 12'h006 ;
		12'hBD0 : douta <= 12'h006 ;
		12'hBD1 : douta <= 12'h006 ;
		12'hBD2 : douta <= 12'h006 ;
		12'hBD3 : douta <= 12'h005 ;
		12'hBD4 : douta <= 12'h005 ;
		12'hBD5 : douta <= 12'h005 ;
		12'hBD6 : douta <= 12'h005 ;
		12'hBD7 : douta <= 12'h005 ;
		12'hBD8 : douta <= 12'h004 ;
		12'hBD9 : douta <= 12'h004 ;
		12'hBDA : douta <= 12'h004 ;
		12'hBDB : douta <= 12'h004 ;
		12'hBDC : douta <= 12'h004 ;
		12'hBDD : douta <= 12'h003 ;
		12'hBDE : douta <= 12'h003 ;
		12'hBDF : douta <= 12'h003 ;
		12'hBE0 : douta <= 12'h003 ;
		12'hBE1 : douta <= 12'h003 ;
		12'hBE2 : douta <= 12'h003 ;
		12'hBE3 : douta <= 12'h003 ;
		12'hBE4 : douta <= 12'h002 ;
		12'hBE5 : douta <= 12'h002 ;
		12'hBE6 : douta <= 12'h002 ;
		12'hBE7 : douta <= 12'h002 ;
		12'hBE8 : douta <= 12'h002 ;
		12'hBE9 : douta <= 12'h002 ;
		12'hBEA : douta <= 12'h002 ;
		12'hBEB : douta <= 12'h002 ;
		12'hBEC : douta <= 12'h001 ;
		12'hBED : douta <= 12'h001 ;
		12'hBEE : douta <= 12'h001 ;
		12'hBEF : douta <= 12'h001 ;
		12'hBF0 : douta <= 12'h001 ;
		12'hBF1 : douta <= 12'h001 ;
		12'hBF2 : douta <= 12'h001 ;
		12'hBF3 : douta <= 12'h001 ;
		12'hBF4 : douta <= 12'h001 ;
		12'hBF5 : douta <= 12'h001 ;
		12'hBF6 : douta <= 12'h001 ;
		12'hBF7 : douta <= 12'h001 ;
		12'hBF8 : douta <= 12'h001 ;
		12'hBF9 : douta <= 12'h001 ;
		12'hBFA : douta <= 12'h001 ;
		12'hBFB : douta <= 12'h001 ;
		12'hBFC : douta <= 12'h001 ;
		12'hBFD : douta <= 12'h001 ;
		12'hBFE : douta <= 12'h001 ;
		12'hBFF : douta <= 12'h001 ;
		12'hC00 : douta <= 12'h000 ;
		12'hC01 : douta <= 12'h001 ;
		12'hC02 : douta <= 12'h001 ;
		12'hC03 : douta <= 12'h001 ;
		12'hC04 : douta <= 12'h001 ;
		12'hC05 : douta <= 12'h001 ;
		12'hC06 : douta <= 12'h001 ;
		12'hC07 : douta <= 12'h001 ;
		12'hC08 : douta <= 12'h001 ;
		12'hC09 : douta <= 12'h001 ;
		12'hC0A : douta <= 12'h001 ;
		12'hC0B : douta <= 12'h001 ;
		12'hC0C : douta <= 12'h001 ;
		12'hC0D : douta <= 12'h001 ;
		12'hC0E : douta <= 12'h001 ;
		12'hC0F : douta <= 12'h001 ;
		12'hC10 : douta <= 12'h001 ;
		12'hC11 : douta <= 12'h001 ;
		12'hC12 : douta <= 12'h001 ;
		12'hC13 : douta <= 12'h001 ;
		12'hC14 : douta <= 12'h001 ;
		12'hC15 : douta <= 12'h002 ;
		12'hC16 : douta <= 12'h002 ;
		12'hC17 : douta <= 12'h002 ;
		12'hC18 : douta <= 12'h002 ;
		12'hC19 : douta <= 12'h002 ;
		12'hC1A : douta <= 12'h002 ;
		12'hC1B : douta <= 12'h002 ;
		12'hC1C : douta <= 12'h002 ;
		12'hC1D : douta <= 12'h003 ;
		12'hC1E : douta <= 12'h003 ;
		12'hC1F : douta <= 12'h003 ;
		12'hC20 : douta <= 12'h003 ;
		12'hC21 : douta <= 12'h003 ;
		12'hC22 : douta <= 12'h003 ;
		12'hC23 : douta <= 12'h003 ;
		12'hC24 : douta <= 12'h004 ;
		12'hC25 : douta <= 12'h004 ;
		12'hC26 : douta <= 12'h004 ;
		12'hC27 : douta <= 12'h004 ;
		12'hC28 : douta <= 12'h004 ;
		12'hC29 : douta <= 12'h005 ;
		12'hC2A : douta <= 12'h005 ;
		12'hC2B : douta <= 12'h005 ;
		12'hC2C : douta <= 12'h005 ;
		12'hC2D : douta <= 12'h005 ;
		12'hC2E : douta <= 12'h006 ;
		12'hC2F : douta <= 12'h006 ;
		12'hC30 : douta <= 12'h006 ;
		12'hC31 : douta <= 12'h006 ;
		12'hC32 : douta <= 12'h007 ;
		12'hC33 : douta <= 12'h007 ;
		12'hC34 : douta <= 12'h007 ;
		12'hC35 : douta <= 12'h007 ;
		12'hC36 : douta <= 12'h008 ;
		12'hC37 : douta <= 12'h008 ;
		12'hC38 : douta <= 12'h008 ;
		12'hC39 : douta <= 12'h008 ;
		12'hC3A : douta <= 12'h009 ;
		12'hC3B : douta <= 12'h009 ;
		12'hC3C : douta <= 12'h009 ;
		12'hC3D : douta <= 12'h009 ;
		12'hC3E : douta <= 12'h00A ;
		12'hC3F : douta <= 12'h00A ;
		12'hC40 : douta <= 12'h00A ;
		12'hC41 : douta <= 12'h00B ;
		12'hC42 : douta <= 12'h00B ;
		12'hC43 : douta <= 12'h00B ;
		12'hC44 : douta <= 12'h00C ;
		12'hC45 : douta <= 12'h00C ;
		12'hC46 : douta <= 12'h00C ;
		12'hC47 : douta <= 12'h00D ;
		12'hC48 : douta <= 12'h00D ;
		12'hC49 : douta <= 12'h00D ;
		12'hC4A : douta <= 12'h00E ;
		12'hC4B : douta <= 12'h00E ;
		12'hC4C : douta <= 12'h00E ;
		12'hC4D : douta <= 12'h00F ;
		12'hC4E : douta <= 12'h00F ;
		12'hC4F : douta <= 12'h010 ;
		12'hC50 : douta <= 12'h010 ;
		12'hC51 : douta <= 12'h010 ;
		12'hC52 : douta <= 12'h011 ;
		12'hC53 : douta <= 12'h011 ;
		12'hC54 : douta <= 12'h011 ;
		12'hC55 : douta <= 12'h012 ;
		12'hC56 : douta <= 12'h012 ;
		12'hC57 : douta <= 12'h013 ;
		12'hC58 : douta <= 12'h013 ;
		12'hC59 : douta <= 12'h014 ;
		12'hC5A : douta <= 12'h014 ;
		12'hC5B : douta <= 12'h014 ;
		12'hC5C : douta <= 12'h015 ;
		12'hC5D : douta <= 12'h015 ;
		12'hC5E : douta <= 12'h016 ;
		12'hC5F : douta <= 12'h016 ;
		12'hC60 : douta <= 12'h017 ;
		12'hC61 : douta <= 12'h017 ;
		12'hC62 : douta <= 12'h018 ;
		12'hC63 : douta <= 12'h018 ;
		12'hC64 : douta <= 12'h019 ;
		12'hC65 : douta <= 12'h019 ;
		12'hC66 : douta <= 12'h01A ;
		12'hC67 : douta <= 12'h01A ;
		12'hC68 : douta <= 12'h01A ;
		12'hC69 : douta <= 12'h01B ;
		12'hC6A : douta <= 12'h01C ;
		12'hC6B : douta <= 12'h01C ;
		12'hC6C : douta <= 12'h01D ;
		12'hC6D : douta <= 12'h01D ;
		12'hC6E : douta <= 12'h01E ;
		12'hC6F : douta <= 12'h01E ;
		12'hC70 : douta <= 12'h01F ;
		12'hC71 : douta <= 12'h01F ;
		12'hC72 : douta <= 12'h020 ;
		12'hC73 : douta <= 12'h020 ;
		12'hC74 : douta <= 12'h021 ;
		12'hC75 : douta <= 12'h021 ;
		12'hC76 : douta <= 12'h022 ;
		12'hC77 : douta <= 12'h023 ;
		12'hC78 : douta <= 12'h023 ;
		12'hC79 : douta <= 12'h024 ;
		12'hC7A : douta <= 12'h024 ;
		12'hC7B : douta <= 12'h025 ;
		12'hC7C : douta <= 12'h025 ;
		12'hC7D : douta <= 12'h026 ;
		12'hC7E : douta <= 12'h027 ;
		12'hC7F : douta <= 12'h027 ;
		12'hC80 : douta <= 12'h028 ;
		12'hC81 : douta <= 12'h028 ;
		12'hC82 : douta <= 12'h029 ;
		12'hC83 : douta <= 12'h02A ;
		12'hC84 : douta <= 12'h02A ;
		12'hC85 : douta <= 12'h02B ;
		12'hC86 : douta <= 12'h02C ;
		12'hC87 : douta <= 12'h02C ;
		12'hC88 : douta <= 12'h02D ;
		12'hC89 : douta <= 12'h02E ;
		12'hC8A : douta <= 12'h02E ;
		12'hC8B : douta <= 12'h02F ;
		12'hC8C : douta <= 12'h030 ;
		12'hC8D : douta <= 12'h030 ;
		12'hC8E : douta <= 12'h031 ;
		12'hC8F : douta <= 12'h032 ;
		12'hC90 : douta <= 12'h032 ;
		12'hC91 : douta <= 12'h033 ;
		12'hC92 : douta <= 12'h034 ;
		12'hC93 : douta <= 12'h034 ;
		12'hC94 : douta <= 12'h035 ;
		12'hC95 : douta <= 12'h036 ;
		12'hC96 : douta <= 12'h036 ;
		12'hC97 : douta <= 12'h037 ;
		12'hC98 : douta <= 12'h038 ;
		12'hC99 : douta <= 12'h039 ;
		12'hC9A : douta <= 12'h039 ;
		12'hC9B : douta <= 12'h03A ;
		12'hC9C : douta <= 12'h03B ;
		12'hC9D : douta <= 12'h03C ;
		12'hC9E : douta <= 12'h03C ;
		12'hC9F : douta <= 12'h03D ;
		12'hCA0 : douta <= 12'h03E ;
		12'hCA1 : douta <= 12'h03F ;
		12'hCA2 : douta <= 12'h03F ;
		12'hCA3 : douta <= 12'h040 ;
		12'hCA4 : douta <= 12'h041 ;
		12'hCA5 : douta <= 12'h042 ;
		12'hCA6 : douta <= 12'h043 ;
		12'hCA7 : douta <= 12'h043 ;
		12'hCA8 : douta <= 12'h044 ;
		12'hCA9 : douta <= 12'h045 ;
		12'hCAA : douta <= 12'h046 ;
		12'hCAB : douta <= 12'h047 ;
		12'hCAC : douta <= 12'h047 ;
		12'hCAD : douta <= 12'h048 ;
		12'hCAE : douta <= 12'h049 ;
		12'hCAF : douta <= 12'h04A ;
		12'hCB0 : douta <= 12'h04B ;
		12'hCB1 : douta <= 12'h04B ;
		12'hCB2 : douta <= 12'h04C ;
		12'hCB3 : douta <= 12'h04D ;
		12'hCB4 : douta <= 12'h04E ;
		12'hCB5 : douta <= 12'h04F ;
		12'hCB6 : douta <= 12'h050 ;
		12'hCB7 : douta <= 12'h051 ;
		12'hCB8 : douta <= 12'h051 ;
		12'hCB9 : douta <= 12'h052 ;
		12'hCBA : douta <= 12'h053 ;
		12'hCBB : douta <= 12'h054 ;
		12'hCBC : douta <= 12'h055 ;
		12'hCBD : douta <= 12'h056 ;
		12'hCBE : douta <= 12'h057 ;
		12'hCBF : douta <= 12'h058 ;
		12'hCC0 : douta <= 12'h059 ;
		12'hCC1 : douta <= 12'h05A ;
		12'hCC2 : douta <= 12'h05A ;
		12'hCC3 : douta <= 12'h05B ;
		12'hCC4 : douta <= 12'h05C ;
		12'hCC5 : douta <= 12'h05D ;
		12'hCC6 : douta <= 12'h05E ;
		12'hCC7 : douta <= 12'h05F ;
		12'hCC8 : douta <= 12'h060 ;
		12'hCC9 : douta <= 12'h061 ;
		12'hCCA : douta <= 12'h062 ;
		12'hCCB : douta <= 12'h063 ;
		12'hCCC : douta <= 12'h064 ;
		12'hCCD : douta <= 12'h065 ;
		12'hCCE : douta <= 12'h066 ;
		12'hCCF : douta <= 12'h067 ;
		12'hCD0 : douta <= 12'h068 ;
		12'hCD1 : douta <= 12'h069 ;
		12'hCD2 : douta <= 12'h06A ;
		12'hCD3 : douta <= 12'h06B ;
		12'hCD4 : douta <= 12'h06C ;
		12'hCD5 : douta <= 12'h06D ;
		12'hCD6 : douta <= 12'h06E ;
		12'hCD7 : douta <= 12'h06F ;
		12'hCD8 : douta <= 12'h070 ;
		12'hCD9 : douta <= 12'h071 ;
		12'hCDA : douta <= 12'h072 ;
		12'hCDB : douta <= 12'h073 ;
		12'hCDC : douta <= 12'h074 ;
		12'hCDD : douta <= 12'h075 ;
		12'hCDE : douta <= 12'h076 ;
		12'hCDF : douta <= 12'h077 ;
		12'hCE0 : douta <= 12'h078 ;
		12'hCE1 : douta <= 12'h079 ;
		12'hCE2 : douta <= 12'h07A ;
		12'hCE3 : douta <= 12'h07B ;
		12'hCE4 : douta <= 12'h07C ;
		12'hCE5 : douta <= 12'h07E ;
		12'hCE6 : douta <= 12'h07F ;
		12'hCE7 : douta <= 12'h080 ;
		12'hCE8 : douta <= 12'h081 ;
		12'hCE9 : douta <= 12'h082 ;
		12'hCEA : douta <= 12'h083 ;
		12'hCEB : douta <= 12'h084 ;
		12'hCEC : douta <= 12'h085 ;
		12'hCED : douta <= 12'h086 ;
		12'hCEE : douta <= 12'h087 ;
		12'hCEF : douta <= 12'h089 ;
		12'hCF0 : douta <= 12'h08A ;
		12'hCF1 : douta <= 12'h08B ;
		12'hCF2 : douta <= 12'h08C ;
		12'hCF3 : douta <= 12'h08D ;
		12'hCF4 : douta <= 12'h08E ;
		12'hCF5 : douta <= 12'h08F ;
		12'hCF6 : douta <= 12'h091 ;
		12'hCF7 : douta <= 12'h092 ;
		12'hCF8 : douta <= 12'h093 ;
		12'hCF9 : douta <= 12'h094 ;
		12'hCFA : douta <= 12'h095 ;
		12'hCFB : douta <= 12'h096 ;
		12'hCFC : douta <= 12'h098 ;
		12'hCFD : douta <= 12'h099 ;
		12'hCFE : douta <= 12'h09A ;
		12'hCFF : douta <= 12'h09B ;
		12'hD00 : douta <= 12'h09C ;
		12'hD01 : douta <= 12'h09E ;
		12'hD02 : douta <= 12'h09F ;
		12'hD03 : douta <= 12'h0A0 ;
		12'hD04 : douta <= 12'h0A1 ;
		12'hD05 : douta <= 12'h0A2 ;
		12'hD06 : douta <= 12'h0A4 ;
		12'hD07 : douta <= 12'h0A5 ;
		12'hD08 : douta <= 12'h0A6 ;
		12'hD09 : douta <= 12'h0A7 ;
		12'hD0A : douta <= 12'h0A9 ;
		12'hD0B : douta <= 12'h0AA ;
		12'hD0C : douta <= 12'h0AB ;
		12'hD0D : douta <= 12'h0AC ;
		12'hD0E : douta <= 12'h0AE ;
		12'hD0F : douta <= 12'h0AF ;
		12'hD10 : douta <= 12'h0B0 ;
		12'hD11 : douta <= 12'h0B1 ;
		12'hD12 : douta <= 12'h0B3 ;
		12'hD13 : douta <= 12'h0B4 ;
		12'hD14 : douta <= 12'h0B5 ;
		12'hD15 : douta <= 12'h0B7 ;
		12'hD16 : douta <= 12'h0B8 ;
		12'hD17 : douta <= 12'h0B9 ;
		12'hD18 : douta <= 12'h0BA ;
		12'hD19 : douta <= 12'h0BC ;
		12'hD1A : douta <= 12'h0BD ;
		12'hD1B : douta <= 12'h0BE ;
		12'hD1C : douta <= 12'h0C0 ;
		12'hD1D : douta <= 12'h0C1 ;
		12'hD1E : douta <= 12'h0C2 ;
		12'hD1F : douta <= 12'h0C4 ;
		12'hD20 : douta <= 12'h0C5 ;
		12'hD21 : douta <= 12'h0C6 ;
		12'hD22 : douta <= 12'h0C8 ;
		12'hD23 : douta <= 12'h0C9 ;
		12'hD24 : douta <= 12'h0CA ;
		12'hD25 : douta <= 12'h0CC ;
		12'hD26 : douta <= 12'h0CD ;
		12'hD27 : douta <= 12'h0CF ;
		12'hD28 : douta <= 12'h0D0 ;
		12'hD29 : douta <= 12'h0D1 ;
		12'hD2A : douta <= 12'h0D3 ;
		12'hD2B : douta <= 12'h0D4 ;
		12'hD2C : douta <= 12'h0D5 ;
		12'hD2D : douta <= 12'h0D7 ;
		12'hD2E : douta <= 12'h0D8 ;
		12'hD2F : douta <= 12'h0DA ;
		12'hD30 : douta <= 12'h0DB ;
		12'hD31 : douta <= 12'h0DC ;
		12'hD32 : douta <= 12'h0DE ;
		12'hD33 : douta <= 12'h0DF ;
		12'hD34 : douta <= 12'h0E1 ;
		12'hD35 : douta <= 12'h0E2 ;
		12'hD36 : douta <= 12'h0E4 ;
		12'hD37 : douta <= 12'h0E5 ;
		12'hD38 : douta <= 12'h0E7 ;
		12'hD39 : douta <= 12'h0E8 ;
		12'hD3A : douta <= 12'h0E9 ;
		12'hD3B : douta <= 12'h0EB ;
		12'hD3C : douta <= 12'h0EC ;
		12'hD3D : douta <= 12'h0EE ;
		12'hD3E : douta <= 12'h0EF ;
		12'hD3F : douta <= 12'h0F1 ;
		12'hD40 : douta <= 12'h0F2 ;
		12'hD41 : douta <= 12'h0F4 ;
		12'hD42 : douta <= 12'h0F5 ;
		12'hD43 : douta <= 12'h0F7 ;
		12'hD44 : douta <= 12'h0F8 ;
		12'hD45 : douta <= 12'h0FA ;
		12'hD46 : douta <= 12'h0FB ;
		12'hD47 : douta <= 12'h0FD ;
		12'hD48 : douta <= 12'h0FE ;
		12'hD49 : douta <= 12'h100 ;
		12'hD4A : douta <= 12'h101 ;
		12'hD4B : douta <= 12'h103 ;
		12'hD4C : douta <= 12'h104 ;
		12'hD4D : douta <= 12'h106 ;
		12'hD4E : douta <= 12'h107 ;
		12'hD4F : douta <= 12'h109 ;
		12'hD50 : douta <= 12'h10A ;
		12'hD51 : douta <= 12'h10C ;
		12'hD52 : douta <= 12'h10E ;
		12'hD53 : douta <= 12'h10F ;
		12'hD54 : douta <= 12'h111 ;
		12'hD55 : douta <= 12'h112 ;
		12'hD56 : douta <= 12'h114 ;
		12'hD57 : douta <= 12'h115 ;
		12'hD58 : douta <= 12'h117 ;
		12'hD59 : douta <= 12'h119 ;
		12'hD5A : douta <= 12'h11A ;
		12'hD5B : douta <= 12'h11C ;
		12'hD5C : douta <= 12'h11D ;
		12'hD5D : douta <= 12'h11F ;
		12'hD5E : douta <= 12'h121 ;
		12'hD5F : douta <= 12'h122 ;
		12'hD60 : douta <= 12'h124 ;
		12'hD61 : douta <= 12'h125 ;
		12'hD62 : douta <= 12'h127 ;
		12'hD63 : douta <= 12'h129 ;
		12'hD64 : douta <= 12'h12A ;
		12'hD65 : douta <= 12'h12C ;
		12'hD66 : douta <= 12'h12D ;
		12'hD67 : douta <= 12'h12F ;
		12'hD68 : douta <= 12'h131 ;
		12'hD69 : douta <= 12'h132 ;
		12'hD6A : douta <= 12'h134 ;
		12'hD6B : douta <= 12'h136 ;
		12'hD6C : douta <= 12'h137 ;
		12'hD6D : douta <= 12'h139 ;
		12'hD6E : douta <= 12'h13B ;
		12'hD6F : douta <= 12'h13C ;
		12'hD70 : douta <= 12'h13E ;
		12'hD71 : douta <= 12'h140 ;
		12'hD72 : douta <= 12'h141 ;
		12'hD73 : douta <= 12'h143 ;
		12'hD74 : douta <= 12'h145 ;
		12'hD75 : douta <= 12'h147 ;
		12'hD76 : douta <= 12'h148 ;
		12'hD77 : douta <= 12'h14A ;
		12'hD78 : douta <= 12'h14C ;
		12'hD79 : douta <= 12'h14D ;
		12'hD7A : douta <= 12'h14F ;
		12'hD7B : douta <= 12'h151 ;
		12'hD7C : douta <= 12'h153 ;
		12'hD7D : douta <= 12'h154 ;
		12'hD7E : douta <= 12'h156 ;
		12'hD7F : douta <= 12'h158 ;
		12'hD80 : douta <= 12'h159 ;
		12'hD81 : douta <= 12'h15B ;
		12'hD82 : douta <= 12'h15D ;
		12'hD83 : douta <= 12'h15F ;
		12'hD84 : douta <= 12'h160 ;
		12'hD85 : douta <= 12'h162 ;
		12'hD86 : douta <= 12'h164 ;
		12'hD87 : douta <= 12'h166 ;
		12'hD88 : douta <= 12'h168 ;
		12'hD89 : douta <= 12'h169 ;
		12'hD8A : douta <= 12'h16B ;
		12'hD8B : douta <= 12'h16D ;
		12'hD8C : douta <= 12'h16F ;
		12'hD8D : douta <= 12'h170 ;
		12'hD8E : douta <= 12'h172 ;
		12'hD8F : douta <= 12'h174 ;
		12'hD90 : douta <= 12'h176 ;
		12'hD91 : douta <= 12'h178 ;
		12'hD92 : douta <= 12'h17A ;
		12'hD93 : douta <= 12'h17B ;
		12'hD94 : douta <= 12'h17D ;
		12'hD95 : douta <= 12'h17F ;
		12'hD96 : douta <= 12'h181 ;
		12'hD97 : douta <= 12'h183 ;
		12'hD98 : douta <= 12'h184 ;
		12'hD99 : douta <= 12'h186 ;
		12'hD9A : douta <= 12'h188 ;
		12'hD9B : douta <= 12'h18A ;
		12'hD9C : douta <= 12'h18C ;
		12'hD9D : douta <= 12'h18E ;
		12'hD9E : douta <= 12'h190 ;
		12'hD9F : douta <= 12'h191 ;
		12'hDA0 : douta <= 12'h193 ;
		12'hDA1 : douta <= 12'h195 ;
		12'hDA2 : douta <= 12'h197 ;
		12'hDA3 : douta <= 12'h199 ;
		12'hDA4 : douta <= 12'h19B ;
		12'hDA5 : douta <= 12'h19D ;
		12'hDA6 : douta <= 12'h19F ;
		12'hDA7 : douta <= 12'h1A1 ;
		12'hDA8 : douta <= 12'h1A2 ;
		12'hDA9 : douta <= 12'h1A4 ;
		12'hDAA : douta <= 12'h1A6 ;
		12'hDAB : douta <= 12'h1A8 ;
		12'hDAC : douta <= 12'h1AA ;
		12'hDAD : douta <= 12'h1AC ;
		12'hDAE : douta <= 12'h1AE ;
		12'hDAF : douta <= 12'h1B0 ;
		12'hDB0 : douta <= 12'h1B2 ;
		12'hDB1 : douta <= 12'h1B4 ;
		12'hDB2 : douta <= 12'h1B6 ;
		12'hDB3 : douta <= 12'h1B8 ;
		12'hDB4 : douta <= 12'h1BA ;
		12'hDB5 : douta <= 12'h1BB ;
		12'hDB6 : douta <= 12'h1BD ;
		12'hDB7 : douta <= 12'h1BF ;
		12'hDB8 : douta <= 12'h1C1 ;
		12'hDB9 : douta <= 12'h1C3 ;
		12'hDBA : douta <= 12'h1C5 ;
		12'hDBB : douta <= 12'h1C7 ;
		12'hDBC : douta <= 12'h1C9 ;
		12'hDBD : douta <= 12'h1CB ;
		12'hDBE : douta <= 12'h1CD ;
		12'hDBF : douta <= 12'h1CF ;
		12'hDC0 : douta <= 12'h1D1 ;
		12'hDC1 : douta <= 12'h1D3 ;
		12'hDC2 : douta <= 12'h1D5 ;
		12'hDC3 : douta <= 12'h1D7 ;
		12'hDC4 : douta <= 12'h1D9 ;
		12'hDC5 : douta <= 12'h1DB ;
		12'hDC6 : douta <= 12'h1DD ;
		12'hDC7 : douta <= 12'h1DF ;
		12'hDC8 : douta <= 12'h1E1 ;
		12'hDC9 : douta <= 12'h1E3 ;
		12'hDCA : douta <= 12'h1E5 ;
		12'hDCB : douta <= 12'h1E7 ;
		12'hDCC : douta <= 12'h1E9 ;
		12'hDCD : douta <= 12'h1EB ;
		12'hDCE : douta <= 12'h1ED ;
		12'hDCF : douta <= 12'h1EF ;
		12'hDD0 : douta <= 12'h1F1 ;
		12'hDD1 : douta <= 12'h1F4 ;
		12'hDD2 : douta <= 12'h1F6 ;
		12'hDD3 : douta <= 12'h1F8 ;
		12'hDD4 : douta <= 12'h1FA ;
		12'hDD5 : douta <= 12'h1FC ;
		12'hDD6 : douta <= 12'h1FE ;
		12'hDD7 : douta <= 12'h200 ;
		12'hDD8 : douta <= 12'h202 ;
		12'hDD9 : douta <= 12'h204 ;
		12'hDDA : douta <= 12'h206 ;
		12'hDDB : douta <= 12'h208 ;
		12'hDDC : douta <= 12'h20A ;
		12'hDDD : douta <= 12'h20C ;
		12'hDDE : douta <= 12'h20F ;
		12'hDDF : douta <= 12'h211 ;
		12'hDE0 : douta <= 12'h213 ;
		12'hDE1 : douta <= 12'h215 ;
		12'hDE2 : douta <= 12'h217 ;
		12'hDE3 : douta <= 12'h219 ;
		12'hDE4 : douta <= 12'h21B ;
		12'hDE5 : douta <= 12'h21D ;
		12'hDE6 : douta <= 12'h21F ;
		12'hDE7 : douta <= 12'h222 ;
		12'hDE8 : douta <= 12'h224 ;
		12'hDE9 : douta <= 12'h226 ;
		12'hDEA : douta <= 12'h228 ;
		12'hDEB : douta <= 12'h22A ;
		12'hDEC : douta <= 12'h22C ;
		12'hDED : douta <= 12'h22E ;
		12'hDEE : douta <= 12'h231 ;
		12'hDEF : douta <= 12'h233 ;
		12'hDF0 : douta <= 12'h235 ;
		12'hDF1 : douta <= 12'h237 ;
		12'hDF2 : douta <= 12'h239 ;
		12'hDF3 : douta <= 12'h23B ;
		12'hDF4 : douta <= 12'h23E ;
		12'hDF5 : douta <= 12'h240 ;
		12'hDF6 : douta <= 12'h242 ;
		12'hDF7 : douta <= 12'h244 ;
		12'hDF8 : douta <= 12'h246 ;
		12'hDF9 : douta <= 12'h249 ;
		12'hDFA : douta <= 12'h24B ;
		12'hDFB : douta <= 12'h24D ;
		12'hDFC : douta <= 12'h24F ;
		12'hDFD : douta <= 12'h251 ;
		12'hDFE : douta <= 12'h254 ;
		12'hDFF : douta <= 12'h256 ;
		12'hE00 : douta <= 12'h258 ;
		12'hE01 : douta <= 12'h25A ;
		12'hE02 : douta <= 12'h25C ;
		12'hE03 : douta <= 12'h25F ;
		12'hE04 : douta <= 12'h261 ;
		12'hE05 : douta <= 12'h263 ;
		12'hE06 : douta <= 12'h265 ;
		12'hE07 : douta <= 12'h268 ;
		12'hE08 : douta <= 12'h26A ;
		12'hE09 : douta <= 12'h26C ;
		12'hE0A : douta <= 12'h26E ;
		12'hE0B : douta <= 12'h271 ;
		12'hE0C : douta <= 12'h273 ;
		12'hE0D : douta <= 12'h275 ;
		12'hE0E : douta <= 12'h277 ;
		12'hE0F : douta <= 12'h27A ;
		12'hE10 : douta <= 12'h27C ;
		12'hE11 : douta <= 12'h27E ;
		12'hE12 : douta <= 12'h281 ;
		12'hE13 : douta <= 12'h283 ;
		12'hE14 : douta <= 12'h285 ;
		12'hE15 : douta <= 12'h287 ;
		12'hE16 : douta <= 12'h28A ;
		12'hE17 : douta <= 12'h28C ;
		12'hE18 : douta <= 12'h28E ;
		12'hE19 : douta <= 12'h291 ;
		12'hE1A : douta <= 12'h293 ;
		12'hE1B : douta <= 12'h295 ;
		12'hE1C : douta <= 12'h298 ;
		12'hE1D : douta <= 12'h29A ;
		12'hE1E : douta <= 12'h29C ;
		12'hE1F : douta <= 12'h29E ;
		12'hE20 : douta <= 12'h2A1 ;
		12'hE21 : douta <= 12'h2A3 ;
		12'hE22 : douta <= 12'h2A5 ;
		12'hE23 : douta <= 12'h2A8 ;
		12'hE24 : douta <= 12'h2AA ;
		12'hE25 : douta <= 12'h2AC ;
		12'hE26 : douta <= 12'h2AF ;
		12'hE27 : douta <= 12'h2B1 ;
		12'hE28 : douta <= 12'h2B4 ;
		12'hE29 : douta <= 12'h2B6 ;
		12'hE2A : douta <= 12'h2B8 ;
		12'hE2B : douta <= 12'h2BB ;
		12'hE2C : douta <= 12'h2BD ;
		12'hE2D : douta <= 12'h2BF ;
		12'hE2E : douta <= 12'h2C2 ;
		12'hE2F : douta <= 12'h2C4 ;
		12'hE30 : douta <= 12'h2C6 ;
		12'hE31 : douta <= 12'h2C9 ;
		12'hE32 : douta <= 12'h2CB ;
		12'hE33 : douta <= 12'h2CE ;
		12'hE34 : douta <= 12'h2D0 ;
		12'hE35 : douta <= 12'h2D2 ;
		12'hE36 : douta <= 12'h2D5 ;
		12'hE37 : douta <= 12'h2D7 ;
		12'hE38 : douta <= 12'h2DA ;
		12'hE39 : douta <= 12'h2DC ;
		12'hE3A : douta <= 12'h2DE ;
		12'hE3B : douta <= 12'h2E1 ;
		12'hE3C : douta <= 12'h2E3 ;
		12'hE3D : douta <= 12'h2E6 ;
		12'hE3E : douta <= 12'h2E8 ;
		12'hE3F : douta <= 12'h2EA ;
		12'hE40 : douta <= 12'h2ED ;
		12'hE41 : douta <= 12'h2EF ;
		12'hE42 : douta <= 12'h2F2 ;
		12'hE43 : douta <= 12'h2F4 ;
		12'hE44 : douta <= 12'h2F7 ;
		12'hE45 : douta <= 12'h2F9 ;
		12'hE46 : douta <= 12'h2FC ;
		12'hE47 : douta <= 12'h2FE ;
		12'hE48 : douta <= 12'h300 ;
		12'hE49 : douta <= 12'h303 ;
		12'hE4A : douta <= 12'h305 ;
		12'hE4B : douta <= 12'h308 ;
		12'hE4C : douta <= 12'h30A ;
		12'hE4D : douta <= 12'h30D ;
		12'hE4E : douta <= 12'h30F ;
		12'hE4F : douta <= 12'h312 ;
		12'hE50 : douta <= 12'h314 ;
		12'hE51 : douta <= 12'h317 ;
		12'hE52 : douta <= 12'h319 ;
		12'hE53 : douta <= 12'h31C ;
		12'hE54 : douta <= 12'h31E ;
		12'hE55 : douta <= 12'h321 ;
		12'hE56 : douta <= 12'h323 ;
		12'hE57 : douta <= 12'h326 ;
		12'hE58 : douta <= 12'h328 ;
		12'hE59 : douta <= 12'h32B ;
		12'hE5A : douta <= 12'h32D ;
		12'hE5B : douta <= 12'h330 ;
		12'hE5C : douta <= 12'h332 ;
		12'hE5D : douta <= 12'h335 ;
		12'hE5E : douta <= 12'h337 ;
		12'hE5F : douta <= 12'h33A ;
		12'hE60 : douta <= 12'h33C ;
		12'hE61 : douta <= 12'h33F ;
		12'hE62 : douta <= 12'h341 ;
		12'hE63 : douta <= 12'h344 ;
		12'hE64 : douta <= 12'h346 ;
		12'hE65 : douta <= 12'h349 ;
		12'hE66 : douta <= 12'h34B ;
		12'hE67 : douta <= 12'h34E ;
		12'hE68 : douta <= 12'h350 ;
		12'hE69 : douta <= 12'h353 ;
		12'hE6A : douta <= 12'h355 ;
		12'hE6B : douta <= 12'h358 ;
		12'hE6C : douta <= 12'h35B ;
		12'hE6D : douta <= 12'h35D ;
		12'hE6E : douta <= 12'h360 ;
		12'hE6F : douta <= 12'h362 ;
		12'hE70 : douta <= 12'h365 ;
		12'hE71 : douta <= 12'h367 ;
		12'hE72 : douta <= 12'h36A ;
		12'hE73 : douta <= 12'h36D ;
		12'hE74 : douta <= 12'h36F ;
		12'hE75 : douta <= 12'h372 ;
		12'hE76 : douta <= 12'h374 ;
		12'hE77 : douta <= 12'h377 ;
		12'hE78 : douta <= 12'h379 ;
		12'hE79 : douta <= 12'h37C ;
		12'hE7A : douta <= 12'h37F ;
		12'hE7B : douta <= 12'h381 ;
		12'hE7C : douta <= 12'h384 ;
		12'hE7D : douta <= 12'h386 ;
		12'hE7E : douta <= 12'h389 ;
		12'hE7F : douta <= 12'h38C ;
		12'hE80 : douta <= 12'h38E ;
		12'hE81 : douta <= 12'h391 ;
		12'hE82 : douta <= 12'h393 ;
		12'hE83 : douta <= 12'h396 ;
		12'hE84 : douta <= 12'h399 ;
		12'hE85 : douta <= 12'h39B ;
		12'hE86 : douta <= 12'h39E ;
		12'hE87 : douta <= 12'h3A1 ;
		12'hE88 : douta <= 12'h3A3 ;
		12'hE89 : douta <= 12'h3A6 ;
		12'hE8A : douta <= 12'h3A8 ;
		12'hE8B : douta <= 12'h3AB ;
		12'hE8C : douta <= 12'h3AE ;
		12'hE8D : douta <= 12'h3B0 ;
		12'hE8E : douta <= 12'h3B3 ;
		12'hE8F : douta <= 12'h3B6 ;
		12'hE90 : douta <= 12'h3B8 ;
		12'hE91 : douta <= 12'h3BB ;
		12'hE92 : douta <= 12'h3BE ;
		12'hE93 : douta <= 12'h3C0 ;
		12'hE94 : douta <= 12'h3C3 ;
		12'hE95 : douta <= 12'h3C6 ;
		12'hE96 : douta <= 12'h3C8 ;
		12'hE97 : douta <= 12'h3CB ;
		12'hE98 : douta <= 12'h3CE ;
		12'hE99 : douta <= 12'h3D0 ;
		12'hE9A : douta <= 12'h3D3 ;
		12'hE9B : douta <= 12'h3D6 ;
		12'hE9C : douta <= 12'h3D8 ;
		12'hE9D : douta <= 12'h3DB ;
		12'hE9E : douta <= 12'h3DE ;
		12'hE9F : douta <= 12'h3E0 ;
		12'hEA0 : douta <= 12'h3E3 ;
		12'hEA1 : douta <= 12'h3E6 ;
		12'hEA2 : douta <= 12'h3E9 ;
		12'hEA3 : douta <= 12'h3EB ;
		12'hEA4 : douta <= 12'h3EE ;
		12'hEA5 : douta <= 12'h3F1 ;
		12'hEA6 : douta <= 12'h3F3 ;
		12'hEA7 : douta <= 12'h3F6 ;
		12'hEA8 : douta <= 12'h3F9 ;
		12'hEA9 : douta <= 12'h3FB ;
		12'hEAA : douta <= 12'h3FE ;
		12'hEAB : douta <= 12'h401 ;
		12'hEAC : douta <= 12'h404 ;
		12'hEAD : douta <= 12'h406 ;
		12'hEAE : douta <= 12'h409 ;
		12'hEAF : douta <= 12'h40C ;
		12'hEB0 : douta <= 12'h40F ;
		12'hEB1 : douta <= 12'h411 ;
		12'hEB2 : douta <= 12'h414 ;
		12'hEB3 : douta <= 12'h417 ;
		12'hEB4 : douta <= 12'h419 ;
		12'hEB5 : douta <= 12'h41C ;
		12'hEB6 : douta <= 12'h41F ;
		12'hEB7 : douta <= 12'h422 ;
		12'hEB8 : douta <= 12'h424 ;
		12'hEB9 : douta <= 12'h427 ;
		12'hEBA : douta <= 12'h42A ;
		12'hEBB : douta <= 12'h42D ;
		12'hEBC : douta <= 12'h42F ;
		12'hEBD : douta <= 12'h432 ;
		12'hEBE : douta <= 12'h435 ;
		12'hEBF : douta <= 12'h438 ;
		12'hEC0 : douta <= 12'h43B ;
		12'hEC1 : douta <= 12'h43D ;
		12'hEC2 : douta <= 12'h440 ;
		12'hEC3 : douta <= 12'h443 ;
		12'hEC4 : douta <= 12'h446 ;
		12'hEC5 : douta <= 12'h448 ;
		12'hEC6 : douta <= 12'h44B ;
		12'hEC7 : douta <= 12'h44E ;
		12'hEC8 : douta <= 12'h451 ;
		12'hEC9 : douta <= 12'h454 ;
		12'hECA : douta <= 12'h456 ;
		12'hECB : douta <= 12'h459 ;
		12'hECC : douta <= 12'h45C ;
		12'hECD : douta <= 12'h45F ;
		12'hECE : douta <= 12'h462 ;
		12'hECF : douta <= 12'h464 ;
		12'hED0 : douta <= 12'h467 ;
		12'hED1 : douta <= 12'h46A ;
		12'hED2 : douta <= 12'h46D ;
		12'hED3 : douta <= 12'h470 ;
		12'hED4 : douta <= 12'h472 ;
		12'hED5 : douta <= 12'h475 ;
		12'hED6 : douta <= 12'h478 ;
		12'hED7 : douta <= 12'h47B ;
		12'hED8 : douta <= 12'h47E ;
		12'hED9 : douta <= 12'h480 ;
		12'hEDA : douta <= 12'h483 ;
		12'hEDB : douta <= 12'h486 ;
		12'hEDC : douta <= 12'h489 ;
		12'hEDD : douta <= 12'h48C ;
		12'hEDE : douta <= 12'h48F ;
		12'hEDF : douta <= 12'h491 ;
		12'hEE0 : douta <= 12'h494 ;
		12'hEE1 : douta <= 12'h497 ;
		12'hEE2 : douta <= 12'h49A ;
		12'hEE3 : douta <= 12'h49D ;
		12'hEE4 : douta <= 12'h4A0 ;
		12'hEE5 : douta <= 12'h4A3 ;
		12'hEE6 : douta <= 12'h4A5 ;
		12'hEE7 : douta <= 12'h4A8 ;
		12'hEE8 : douta <= 12'h4AB ;
		12'hEE9 : douta <= 12'h4AE ;
		12'hEEA : douta <= 12'h4B1 ;
		12'hEEB : douta <= 12'h4B4 ;
		12'hEEC : douta <= 12'h4B7 ;
		12'hEED : douta <= 12'h4B9 ;
		12'hEEE : douta <= 12'h4BC ;
		12'hEEF : douta <= 12'h4BF ;
		12'hEF0 : douta <= 12'h4C2 ;
		12'hEF1 : douta <= 12'h4C5 ;
		12'hEF2 : douta <= 12'h4C8 ;
		12'hEF3 : douta <= 12'h4CB ;
		12'hEF4 : douta <= 12'h4CD ;
		12'hEF5 : douta <= 12'h4D0 ;
		12'hEF6 : douta <= 12'h4D3 ;
		12'hEF7 : douta <= 12'h4D6 ;
		12'hEF8 : douta <= 12'h4D9 ;
		12'hEF9 : douta <= 12'h4DC ;
		12'hEFA : douta <= 12'h4DF ;
		12'hEFB : douta <= 12'h4E2 ;
		12'hEFC : douta <= 12'h4E5 ;
		12'hEFD : douta <= 12'h4E7 ;
		12'hEFE : douta <= 12'h4EA ;
		12'hEFF : douta <= 12'h4ED ;
		12'hF00 : douta <= 12'h4F0 ;
		12'hF01 : douta <= 12'h4F3 ;
		12'hF02 : douta <= 12'h4F6 ;
		12'hF03 : douta <= 12'h4F9 ;
		12'hF04 : douta <= 12'h4FC ;
		12'hF05 : douta <= 12'h4FF ;
		12'hF06 : douta <= 12'h502 ;
		12'hF07 : douta <= 12'h504 ;
		12'hF08 : douta <= 12'h507 ;
		12'hF09 : douta <= 12'h50A ;
		12'hF0A : douta <= 12'h50D ;
		12'hF0B : douta <= 12'h510 ;
		12'hF0C : douta <= 12'h513 ;
		12'hF0D : douta <= 12'h516 ;
		12'hF0E : douta <= 12'h519 ;
		12'hF0F : douta <= 12'h51C ;
		12'hF10 : douta <= 12'h51F ;
		12'hF11 : douta <= 12'h522 ;
		12'hF12 : douta <= 12'h525 ;
		12'hF13 : douta <= 12'h528 ;
		12'hF14 : douta <= 12'h52B ;
		12'hF15 : douta <= 12'h52D ;
		12'hF16 : douta <= 12'h530 ;
		12'hF17 : douta <= 12'h533 ;
		12'hF18 : douta <= 12'h536 ;
		12'hF19 : douta <= 12'h539 ;
		12'hF1A : douta <= 12'h53C ;
		12'hF1B : douta <= 12'h53F ;
		12'hF1C : douta <= 12'h542 ;
		12'hF1D : douta <= 12'h545 ;
		12'hF1E : douta <= 12'h548 ;
		12'hF1F : douta <= 12'h54B ;
		12'hF20 : douta <= 12'h54E ;
		12'hF21 : douta <= 12'h551 ;
		12'hF22 : douta <= 12'h554 ;
		12'hF23 : douta <= 12'h557 ;
		12'hF24 : douta <= 12'h55A ;
		12'hF25 : douta <= 12'h55D ;
		12'hF26 : douta <= 12'h560 ;
		12'hF27 : douta <= 12'h563 ;
		12'hF28 : douta <= 12'h566 ;
		12'hF29 : douta <= 12'h569 ;
		12'hF2A : douta <= 12'h56C ;
		12'hF2B : douta <= 12'h56F ;
		12'hF2C : douta <= 12'h571 ;
		12'hF2D : douta <= 12'h574 ;
		12'hF2E : douta <= 12'h577 ;
		12'hF2F : douta <= 12'h57A ;
		12'hF30 : douta <= 12'h57D ;
		12'hF31 : douta <= 12'h580 ;
		12'hF32 : douta <= 12'h583 ;
		12'hF33 : douta <= 12'h586 ;
		12'hF34 : douta <= 12'h589 ;
		12'hF35 : douta <= 12'h58C ;
		12'hF36 : douta <= 12'h58F ;
		12'hF37 : douta <= 12'h592 ;
		12'hF38 : douta <= 12'h595 ;
		12'hF39 : douta <= 12'h598 ;
		12'hF3A : douta <= 12'h59B ;
		12'hF3B : douta <= 12'h59E ;
		12'hF3C : douta <= 12'h5A1 ;
		12'hF3D : douta <= 12'h5A4 ;
		12'hF3E : douta <= 12'h5A7 ;
		12'hF3F : douta <= 12'h5AA ;
		12'hF40 : douta <= 12'h5AD ;
		12'hF41 : douta <= 12'h5B0 ;
		12'hF42 : douta <= 12'h5B3 ;
		12'hF43 : douta <= 12'h5B6 ;
		12'hF44 : douta <= 12'h5B9 ;
		12'hF45 : douta <= 12'h5BC ;
		12'hF46 : douta <= 12'h5BF ;
		12'hF47 : douta <= 12'h5C2 ;
		12'hF48 : douta <= 12'h5C5 ;
		12'hF49 : douta <= 12'h5C8 ;
		12'hF4A : douta <= 12'h5CB ;
		12'hF4B : douta <= 12'h5CE ;
		12'hF4C : douta <= 12'h5D1 ;
		12'hF4D : douta <= 12'h5D4 ;
		12'hF4E : douta <= 12'h5D7 ;
		12'hF4F : douta <= 12'h5DB ;
		12'hF50 : douta <= 12'h5DE ;
		12'hF51 : douta <= 12'h5E1 ;
		12'hF52 : douta <= 12'h5E4 ;
		12'hF53 : douta <= 12'h5E7 ;
		12'hF54 : douta <= 12'h5EA ;
		12'hF55 : douta <= 12'h5ED ;
		12'hF56 : douta <= 12'h5F0 ;
		12'hF57 : douta <= 12'h5F3 ;
		12'hF58 : douta <= 12'h5F6 ;
		12'hF59 : douta <= 12'h5F9 ;
		12'hF5A : douta <= 12'h5FC ;
		12'hF5B : douta <= 12'h5FF ;
		12'hF5C : douta <= 12'h602 ;
		12'hF5D : douta <= 12'h605 ;
		12'hF5E : douta <= 12'h608 ;
		12'hF5F : douta <= 12'h60B ;
		12'hF60 : douta <= 12'h60E ;
		12'hF61 : douta <= 12'h611 ;
		12'hF62 : douta <= 12'h614 ;
		12'hF63 : douta <= 12'h617 ;
		12'hF64 : douta <= 12'h61A ;
		12'hF65 : douta <= 12'h61D ;
		12'hF66 : douta <= 12'h620 ;
		12'hF67 : douta <= 12'h623 ;
		12'hF68 : douta <= 12'h627 ;
		12'hF69 : douta <= 12'h62A ;
		12'hF6A : douta <= 12'h62D ;
		12'hF6B : douta <= 12'h630 ;
		12'hF6C : douta <= 12'h633 ;
		12'hF6D : douta <= 12'h636 ;
		12'hF6E : douta <= 12'h639 ;
		12'hF6F : douta <= 12'h63C ;
		12'hF70 : douta <= 12'h63F ;
		12'hF71 : douta <= 12'h642 ;
		12'hF72 : douta <= 12'h645 ;
		12'hF73 : douta <= 12'h648 ;
		12'hF74 : douta <= 12'h64B ;
		12'hF75 : douta <= 12'h64E ;
		12'hF76 : douta <= 12'h651 ;
		12'hF77 : douta <= 12'h654 ;
		12'hF78 : douta <= 12'h658 ;
		12'hF79 : douta <= 12'h65B ;
		12'hF7A : douta <= 12'h65E ;
		12'hF7B : douta <= 12'h661 ;
		12'hF7C : douta <= 12'h664 ;
		12'hF7D : douta <= 12'h667 ;
		12'hF7E : douta <= 12'h66A ;
		12'hF7F : douta <= 12'h66D ;
		12'hF80 : douta <= 12'h670 ;
		12'hF81 : douta <= 12'h673 ;
		12'hF82 : douta <= 12'h676 ;
		12'hF83 : douta <= 12'h679 ;
		12'hF84 : douta <= 12'h67C ;
		12'hF85 : douta <= 12'h680 ;
		12'hF86 : douta <= 12'h683 ;
		12'hF87 : douta <= 12'h686 ;
		12'hF88 : douta <= 12'h689 ;
		12'hF89 : douta <= 12'h68C ;
		12'hF8A : douta <= 12'h68F ;
		12'hF8B : douta <= 12'h692 ;
		12'hF8C : douta <= 12'h695 ;
		12'hF8D : douta <= 12'h698 ;
		12'hF8E : douta <= 12'h69B ;
		12'hF8F : douta <= 12'h69E ;
		12'hF90 : douta <= 12'h6A2 ;
		12'hF91 : douta <= 12'h6A5 ;
		12'hF92 : douta <= 12'h6A8 ;
		12'hF93 : douta <= 12'h6AB ;
		12'hF94 : douta <= 12'h6AE ;
		12'hF95 : douta <= 12'h6B1 ;
		12'hF96 : douta <= 12'h6B4 ;
		12'hF97 : douta <= 12'h6B7 ;
		12'hF98 : douta <= 12'h6BA ;
		12'hF99 : douta <= 12'h6BD ;
		12'hF9A : douta <= 12'h6C1 ;
		12'hF9B : douta <= 12'h6C4 ;
		12'hF9C : douta <= 12'h6C7 ;
		12'hF9D : douta <= 12'h6CA ;
		12'hF9E : douta <= 12'h6CD ;
		12'hF9F : douta <= 12'h6D0 ;
		12'hFA0 : douta <= 12'h6D3 ;
		12'hFA1 : douta <= 12'h6D6 ;
		12'hFA2 : douta <= 12'h6D9 ;
		12'hFA3 : douta <= 12'h6DC ;
		12'hFA4 : douta <= 12'h6E0 ;
		12'hFA5 : douta <= 12'h6E3 ;
		12'hFA6 : douta <= 12'h6E6 ;
		12'hFA7 : douta <= 12'h6E9 ;
		12'hFA8 : douta <= 12'h6EC ;
		12'hFA9 : douta <= 12'h6EF ;
		12'hFAA : douta <= 12'h6F2 ;
		12'hFAB : douta <= 12'h6F5 ;
		12'hFAC : douta <= 12'h6F8 ;
		12'hFAD : douta <= 12'h6FC ;
		12'hFAE : douta <= 12'h6FF ;
		12'hFAF : douta <= 12'h702 ;
		12'hFB0 : douta <= 12'h705 ;
		12'hFB1 : douta <= 12'h708 ;
		12'hFB2 : douta <= 12'h70B ;
		12'hFB3 : douta <= 12'h70E ;
		12'hFB4 : douta <= 12'h711 ;
		12'hFB5 : douta <= 12'h715 ;
		12'hFB6 : douta <= 12'h718 ;
		12'hFB7 : douta <= 12'h71B ;
		12'hFB8 : douta <= 12'h71E ;
		12'hFB9 : douta <= 12'h721 ;
		12'hFBA : douta <= 12'h724 ;
		12'hFBB : douta <= 12'h727 ;
		12'hFBC : douta <= 12'h72A ;
		12'hFBD : douta <= 12'h72D ;
		12'hFBE : douta <= 12'h731 ;
		12'hFBF : douta <= 12'h734 ;
		12'hFC0 : douta <= 12'h737 ;
		12'hFC1 : douta <= 12'h73A ;
		12'hFC2 : douta <= 12'h73D ;
		12'hFC3 : douta <= 12'h740 ;
		12'hFC4 : douta <= 12'h743 ;
		12'hFC5 : douta <= 12'h746 ;
		12'hFC6 : douta <= 12'h74A ;
		12'hFC7 : douta <= 12'h74D ;
		12'hFC8 : douta <= 12'h750 ;
		12'hFC9 : douta <= 12'h753 ;
		12'hFCA : douta <= 12'h756 ;
		12'hFCB : douta <= 12'h759 ;
		12'hFCC : douta <= 12'h75C ;
		12'hFCD : douta <= 12'h760 ;
		12'hFCE : douta <= 12'h763 ;
		12'hFCF : douta <= 12'h766 ;
		12'hFD0 : douta <= 12'h769 ;
		12'hFD1 : douta <= 12'h76C ;
		12'hFD2 : douta <= 12'h76F ;
		12'hFD3 : douta <= 12'h772 ;
		12'hFD4 : douta <= 12'h775 ;
		12'hFD5 : douta <= 12'h779 ;
		12'hFD6 : douta <= 12'h77C ;
		12'hFD7 : douta <= 12'h77F ;
		12'hFD8 : douta <= 12'h782 ;
		12'hFD9 : douta <= 12'h785 ;
		12'hFDA : douta <= 12'h788 ;
		12'hFDB : douta <= 12'h78B ;
		12'hFDC : douta <= 12'h78F ;
		12'hFDD : douta <= 12'h792 ;
		12'hFDE : douta <= 12'h795 ;
		12'hFDF : douta <= 12'h798 ;
		12'hFE0 : douta <= 12'h79B ;
		12'hFE1 : douta <= 12'h79E ;
		12'hFE2 : douta <= 12'h7A1 ;
		12'hFE3 : douta <= 12'h7A4 ;
		12'hFE4 : douta <= 12'h7A8 ;
		12'hFE5 : douta <= 12'h7AB ;
		12'hFE6 : douta <= 12'h7AE ;
		12'hFE7 : douta <= 12'h7B1 ;
		12'hFE8 : douta <= 12'h7B4 ;
		12'hFE9 : douta <= 12'h7B7 ;
		12'hFEA : douta <= 12'h7BA ;
		12'hFEB : douta <= 12'h7BE ;
		12'hFEC : douta <= 12'h7C1 ;
		12'hFED : douta <= 12'h7C4 ;
		12'hFEE : douta <= 12'h7C7 ;
		12'hFEF : douta <= 12'h7CA ;
		12'hFF0 : douta <= 12'h7CD ;
		12'hFF1 : douta <= 12'h7D0 ;
		12'hFF2 : douta <= 12'h7D4 ;
		12'hFF3 : douta <= 12'h7D7 ;
		12'hFF4 : douta <= 12'h7DA ;
		12'hFF5 : douta <= 12'h7DD ;
		12'hFF6 : douta <= 12'h7E0 ;
		12'hFF7 : douta <= 12'h7E3 ;
		12'hFF8 : douta <= 12'h7E6 ;
		12'hFF9 : douta <= 12'h7EA ;
		12'hFFA : douta <= 12'h7ED ;
		12'hFFB : douta <= 12'h7F0 ;
		12'hFFC : douta <= 12'h7F3 ;
		12'hFFD : douta <= 12'h7F6 ;
		12'hFFE : douta <= 12'h7F9 ;
		12'hFFF : douta <= 12'h7FC ;
		endcase
end	

endmodule