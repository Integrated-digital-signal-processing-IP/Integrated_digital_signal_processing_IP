module usin_rom
(
input	wire			clk		,
input	wire			rst 	,
input	wire	[11:0]	addr	,
output	reg 	[11:0]	dout
);
		
always@ (posedge clk, negedge rst)
begin
	if (!rst)
		dout <= 0;
	else
		case ( addra )
		12'h000 : dout <= 12'h800;
		12'h001 : dout <= 12'h803;
		12'h002 : dout <= 12'h806;
		12'h003 : dout <= 12'h809;
		12'h004 : dout <= 12'h80C;
		12'h005 : dout <= 12'h80F;
		12'h006 : dout <= 12'h812;
		12'h007 : dout <= 12'h815;
		12'h008 : dout <= 12'h819;
		12'h009 : dout <= 12'h81C;
		12'h00A : dout <= 12'h81F;
		12'h00B : dout <= 12'h822;
		12'h00C : dout <= 12'h825;
		12'h00D : dout <= 12'h828;
		12'h00E : dout <= 12'h82B;
		12'h00F : dout <= 12'h82F;
		12'h010 : dout <= 12'h832;
		12'h011 : dout <= 12'h835;
		12'h012 : dout <= 12'h838;
		12'h013 : dout <= 12'h83B;
		12'h014 : dout <= 12'h83E;
		12'h015 : dout <= 12'h841;
		12'h016 : dout <= 12'h845;
		12'h017 : dout <= 12'h848;
		12'h018 : dout <= 12'h84B;
		12'h019 : dout <= 12'h84E;
		12'h01A : dout <= 12'h851;
		12'h01B : dout <= 12'h854;
		12'h01C : dout <= 12'h857;
		12'h01D : dout <= 12'h85B;
		12'h01E : dout <= 12'h85E;
		12'h01F : dout <= 12'h861;
		12'h020 : dout <= 12'h864;
		12'h021 : dout <= 12'h867;
		12'h022 : dout <= 12'h86A;
		12'h023 : dout <= 12'h86D;
		12'h024 : dout <= 12'h870;
		12'h025 : dout <= 12'h874;
		12'h026 : dout <= 12'h877;
		12'h027 : dout <= 12'h87A;
		12'h028 : dout <= 12'h87D;
		12'h029 : dout <= 12'h880;
		12'h02A : dout <= 12'h883;
		12'h02B : dout <= 12'h886;
		12'h02C : dout <= 12'h88A;
		12'h02D : dout <= 12'h88D;
		12'h02E : dout <= 12'h890;
		12'h02F : dout <= 12'h893;
		12'h030 : dout <= 12'h896;
		12'h031 : dout <= 12'h899;
		12'h032 : dout <= 12'h89C;
		12'h033 : dout <= 12'h89F;
		12'h034 : dout <= 12'h8A3;
		12'h035 : dout <= 12'h8A6;
		12'h036 : dout <= 12'h8A9;
		12'h037 : dout <= 12'h8AC;
		12'h038 : dout <= 12'h8AF;
		12'h039 : dout <= 12'h8B2;
		12'h03A : dout <= 12'h8B5;
		12'h03B : dout <= 12'h8B9;
		12'h03C : dout <= 12'h8BC;
		12'h03D : dout <= 12'h8BF;
		12'h03E : dout <= 12'h8C2;
		12'h03F : dout <= 12'h8C5;
		12'h040 : dout <= 12'h8C8;
		12'h041 : dout <= 12'h8CB;
		12'h042 : dout <= 12'h8CE;
		12'h043 : dout <= 12'h8D2;
		12'h044 : dout <= 12'h8D5;
		12'h045 : dout <= 12'h8D8;
		12'h046 : dout <= 12'h8DB;
		12'h047 : dout <= 12'h8DE;
		12'h048 : dout <= 12'h8E1;
		12'h049 : dout <= 12'h8E4;
		12'h04A : dout <= 12'h8E7;
		12'h04B : dout <= 12'h8EA;
		12'h04C : dout <= 12'h8EE;
		12'h04D : dout <= 12'h8F1;
		12'h04E : dout <= 12'h8F4;
		12'h04F : dout <= 12'h8F7;
		12'h050 : dout <= 12'h8FA;
		12'h051 : dout <= 12'h8FD;
		12'h052 : dout <= 12'h900;
		12'h053 : dout <= 12'h903;
		12'h054 : dout <= 12'h907;
		12'h055 : dout <= 12'h90A;
		12'h056 : dout <= 12'h90D;
		12'h057 : dout <= 12'h910;
		12'h058 : dout <= 12'h913;
		12'h059 : dout <= 12'h916;
		12'h05A : dout <= 12'h919;
		12'h05B : dout <= 12'h91C;
		12'h05C : dout <= 12'h91F;
		12'h05D : dout <= 12'h923;
		12'h05E : dout <= 12'h926;
		12'h05F : dout <= 12'h929;
		12'h060 : dout <= 12'h92C;
		12'h061 : dout <= 12'h92F;
		12'h062 : dout <= 12'h932;
		12'h063 : dout <= 12'h935;
		12'h064 : dout <= 12'h938;
		12'h065 : dout <= 12'h93B;
		12'h066 : dout <= 12'h93E;
		12'h067 : dout <= 12'h942;
		12'h068 : dout <= 12'h945;
		12'h069 : dout <= 12'h948;
		12'h06A : dout <= 12'h94B;
		12'h06B : dout <= 12'h94E;
		12'h06C : dout <= 12'h951;
		12'h06D : dout <= 12'h954;
		12'h06E : dout <= 12'h957;
		12'h06F : dout <= 12'h95A;
		12'h070 : dout <= 12'h95D;
		12'h071 : dout <= 12'h961;
		12'h072 : dout <= 12'h964;
		12'h073 : dout <= 12'h967;
		12'h074 : dout <= 12'h96A;
		12'h075 : dout <= 12'h96D;
		12'h076 : dout <= 12'h970;
		12'h077 : dout <= 12'h973;
		12'h078 : dout <= 12'h976;
		12'h079 : dout <= 12'h979;
		12'h07A : dout <= 12'h97C;
		12'h07B : dout <= 12'h97F;
		12'h07C : dout <= 12'h983;
		12'h07D : dout <= 12'h986;
		12'h07E : dout <= 12'h989;
		12'h07F : dout <= 12'h98C;
		12'h080 : dout <= 12'h98F;
		12'h081 : dout <= 12'h992;
		12'h082 : dout <= 12'h995;
		12'h083 : dout <= 12'h998;
		12'h084 : dout <= 12'h99B;
		12'h085 : dout <= 12'h99E;
		12'h086 : dout <= 12'h9A1;
		12'h087 : dout <= 12'h9A4;
		12'h088 : dout <= 12'h9A7;
		12'h089 : dout <= 12'h9AB;
		12'h08A : dout <= 12'h9AE;
		12'h08B : dout <= 12'h9B1;
		12'h08C : dout <= 12'h9B4;
		12'h08D : dout <= 12'h9B7;
		12'h08E : dout <= 12'h9BA;
		12'h08F : dout <= 12'h9BD;
		12'h090 : dout <= 12'h9C0;
		12'h091 : dout <= 12'h9C3;
		12'h092 : dout <= 12'h9C6;
		12'h093 : dout <= 12'h9C9;
		12'h094 : dout <= 12'h9CC;
		12'h095 : dout <= 12'h9CF;
		12'h096 : dout <= 12'h9D2;
		12'h097 : dout <= 12'h9D5;
		12'h098 : dout <= 12'h9D8;
		12'h099 : dout <= 12'h9DC;
		12'h09A : dout <= 12'h9DF;
		12'h09B : dout <= 12'h9E2;
		12'h09C : dout <= 12'h9E5;
		12'h09D : dout <= 12'h9E8;
		12'h09E : dout <= 12'h9EB;
		12'h09F : dout <= 12'h9EE;
		12'h0A0 : dout <= 12'h9F1;
		12'h0A1 : dout <= 12'h9F4;
		12'h0A2 : dout <= 12'h9F7;
		12'h0A3 : dout <= 12'h9FA;
		12'h0A4 : dout <= 12'h9FD;
		12'h0A5 : dout <= 12'hA00;
		12'h0A6 : dout <= 12'hA03;
		12'h0A7 : dout <= 12'hA06;
		12'h0A8 : dout <= 12'hA09;
		12'h0A9 : dout <= 12'hA0C;
		12'h0AA : dout <= 12'hA0F;
		12'h0AB : dout <= 12'hA12;
		12'h0AC : dout <= 12'hA15;
		12'h0AD : dout <= 12'hA18;
		12'h0AE : dout <= 12'hA1B;
		12'h0AF : dout <= 12'hA1E;
		12'h0B0 : dout <= 12'hA21;
		12'h0B1 : dout <= 12'hA24;
		12'h0B2 : dout <= 12'hA28;
		12'h0B3 : dout <= 12'hA2B;
		12'h0B4 : dout <= 12'hA2E;
		12'h0B5 : dout <= 12'hA31;
		12'h0B6 : dout <= 12'hA34;
		12'h0B7 : dout <= 12'hA37;
		12'h0B8 : dout <= 12'hA3A;
		12'h0B9 : dout <= 12'hA3D;
		12'h0BA : dout <= 12'hA40;
		12'h0BB : dout <= 12'hA43;
		12'h0BC : dout <= 12'hA46;
		12'h0BD : dout <= 12'hA49;
		12'h0BE : dout <= 12'hA4C;
		12'h0BF : dout <= 12'hA4F;
		12'h0C0 : dout <= 12'hA52;
		12'h0C1 : dout <= 12'hA55;
		12'h0C2 : dout <= 12'hA58;
		12'h0C3 : dout <= 12'hA5B;
		12'h0C4 : dout <= 12'hA5E;
		12'h0C5 : dout <= 12'hA61;
		12'h0C6 : dout <= 12'hA64;
		12'h0C7 : dout <= 12'hA67;
		12'h0C8 : dout <= 12'hA6A;
		12'h0C9 : dout <= 12'hA6D;
		12'h0CA : dout <= 12'hA70;
		12'h0CB : dout <= 12'hA73;
		12'h0CC : dout <= 12'hA76;
		12'h0CD : dout <= 12'hA79;
		12'h0CE : dout <= 12'hA7C;
		12'h0CF : dout <= 12'hA7F;
		12'h0D0 : dout <= 12'hA82;
		12'h0D1 : dout <= 12'hA85;
		12'h0D2 : dout <= 12'hA88;
		12'h0D3 : dout <= 12'hA8B;
		12'h0D4 : dout <= 12'hA8E;
		12'h0D5 : dout <= 12'hA90;
		12'h0D6 : dout <= 12'hA93;
		12'h0D7 : dout <= 12'hA96;
		12'h0D8 : dout <= 12'hA99;
		12'h0D9 : dout <= 12'hA9C;
		12'h0DA : dout <= 12'hA9F;
		12'h0DB : dout <= 12'hAA2;
		12'h0DC : dout <= 12'hAA5;
		12'h0DD : dout <= 12'hAA8;
		12'h0DE : dout <= 12'hAAB;
		12'h0DF : dout <= 12'hAAE;
		12'h0E0 : dout <= 12'hAB1;
		12'h0E1 : dout <= 12'hAB4;
		12'h0E2 : dout <= 12'hAB7;
		12'h0E3 : dout <= 12'hABA;
		12'h0E4 : dout <= 12'hABD;
		12'h0E5 : dout <= 12'hAC0;
		12'h0E6 : dout <= 12'hAC3;
		12'h0E7 : dout <= 12'hAC6;
		12'h0E8 : dout <= 12'hAC9;
		12'h0E9 : dout <= 12'hACC;
		12'h0EA : dout <= 12'hACF;
		12'h0EB : dout <= 12'hAD2;
		12'h0EC : dout <= 12'hAD4;
		12'h0ED : dout <= 12'hAD7;
		12'h0EE : dout <= 12'hADA;
		12'h0EF : dout <= 12'hADD;
		12'h0F0 : dout <= 12'hAE0;
		12'h0F1 : dout <= 12'hAE3;
		12'h0F2 : dout <= 12'hAE6;
		12'h0F3 : dout <= 12'hAE9;
		12'h0F4 : dout <= 12'hAEC;
		12'h0F5 : dout <= 12'hAEF;
		12'h0F6 : dout <= 12'hAF2;
		12'h0F7 : dout <= 12'hAF5;
		12'h0F8 : dout <= 12'hAF8;
		12'h0F9 : dout <= 12'hAFB;
		12'h0FA : dout <= 12'hAFD;
		12'h0FB : dout <= 12'hB00;
		12'h0FC : dout <= 12'hB03;
		12'h0FD : dout <= 12'hB06;
		12'h0FE : dout <= 12'hB09;
		12'h0FF : dout <= 12'hB0C;
		12'h100 : dout <= 12'hB0F;
		12'h101 : dout <= 12'hB12;
		12'h102 : dout <= 12'hB15;
		12'h103 : dout <= 12'hB18;
		12'h104 : dout <= 12'hB1A;
		12'h105 : dout <= 12'hB1D;
		12'h106 : dout <= 12'hB20;
		12'h107 : dout <= 12'hB23;
		12'h108 : dout <= 12'hB26;
		12'h109 : dout <= 12'hB29;
		12'h10A : dout <= 12'hB2C;
		12'h10B : dout <= 12'hB2F;
		12'h10C : dout <= 12'hB32;
		12'h10D : dout <= 12'hB34;
		12'h10E : dout <= 12'hB37;
		12'h10F : dout <= 12'hB3A;
		12'h110 : dout <= 12'hB3D;
		12'h111 : dout <= 12'hB40;
		12'h112 : dout <= 12'hB43;
		12'h113 : dout <= 12'hB46;
		12'h114 : dout <= 12'hB48;
		12'h115 : dout <= 12'hB4B;
		12'h116 : dout <= 12'hB4E;
		12'h117 : dout <= 12'hB51;
		12'h118 : dout <= 12'hB54;
		12'h119 : dout <= 12'hB57;
		12'h11A : dout <= 12'hB5A;
		12'h11B : dout <= 12'hB5C;
		12'h11C : dout <= 12'hB5F;
		12'h11D : dout <= 12'hB62;
		12'h11E : dout <= 12'hB65;
		12'h11F : dout <= 12'hB68;
		12'h120 : dout <= 12'hB6B;
		12'h121 : dout <= 12'hB6E;
		12'h122 : dout <= 12'hB70;
		12'h123 : dout <= 12'hB73;
		12'h124 : dout <= 12'hB76;
		12'h125 : dout <= 12'hB79;
		12'h126 : dout <= 12'hB7C;
		12'h127 : dout <= 12'hB7F;
		12'h128 : dout <= 12'hB81;
		12'h129 : dout <= 12'hB84;
		12'h12A : dout <= 12'hB87;
		12'h12B : dout <= 12'hB8A;
		12'h12C : dout <= 12'hB8D;
		12'h12D : dout <= 12'hB8F;
		12'h12E : dout <= 12'hB92;
		12'h12F : dout <= 12'hB95;
		12'h130 : dout <= 12'hB98;
		12'h131 : dout <= 12'hB9B;
		12'h132 : dout <= 12'hB9D;
		12'h133 : dout <= 12'hBA0;
		12'h134 : dout <= 12'hBA3;
		12'h135 : dout <= 12'hBA6;
		12'h136 : dout <= 12'hBA9;
		12'h137 : dout <= 12'hBAB;
		12'h138 : dout <= 12'hBAE;
		12'h139 : dout <= 12'hBB1;
		12'h13A : dout <= 12'hBB4;
		12'h13B : dout <= 12'hBB7;
		12'h13C : dout <= 12'hBB9;
		12'h13D : dout <= 12'hBBC;
		12'h13E : dout <= 12'hBBF;
		12'h13F : dout <= 12'hBC2;
		12'h140 : dout <= 12'hBC4;
		12'h141 : dout <= 12'hBC7;
		12'h142 : dout <= 12'hBCA;
		12'h143 : dout <= 12'hBCD;
		12'h144 : dout <= 12'hBD0;
		12'h145 : dout <= 12'hBD2;
		12'h146 : dout <= 12'hBD5;
		12'h147 : dout <= 12'hBD8;
		12'h148 : dout <= 12'hBDB;
		12'h149 : dout <= 12'hBDD;
		12'h14A : dout <= 12'hBE0;
		12'h14B : dout <= 12'hBE3;
		12'h14C : dout <= 12'hBE6;
		12'h14D : dout <= 12'hBE8;
		12'h14E : dout <= 12'hBEB;
		12'h14F : dout <= 12'hBEE;
		12'h150 : dout <= 12'hBF0;
		12'h151 : dout <= 12'hBF3;
		12'h152 : dout <= 12'hBF6;
		12'h153 : dout <= 12'hBF9;
		12'h154 : dout <= 12'hBFB;
		12'h155 : dout <= 12'hBFE;
		12'h156 : dout <= 12'hC01;
		12'h157 : dout <= 12'hC04;
		12'h158 : dout <= 12'hC06;
		12'h159 : dout <= 12'hC09;
		12'h15A : dout <= 12'hC0C;
		12'h15B : dout <= 12'hC0E;
		12'h15C : dout <= 12'hC11;
		12'h15D : dout <= 12'hC14;
		12'h15E : dout <= 12'hC16;
		12'h15F : dout <= 12'hC19;
		12'h160 : dout <= 12'hC1C;
		12'h161 : dout <= 12'hC1F;
		12'h162 : dout <= 12'hC21;
		12'h163 : dout <= 12'hC24;
		12'h164 : dout <= 12'hC27;
		12'h165 : dout <= 12'hC29;
		12'h166 : dout <= 12'hC2C;
		12'h167 : dout <= 12'hC2F;
		12'h168 : dout <= 12'hC31;
		12'h169 : dout <= 12'hC34;
		12'h16A : dout <= 12'hC37;
		12'h16B : dout <= 12'hC39;
		12'h16C : dout <= 12'hC3C;
		12'h16D : dout <= 12'hC3F;
		12'h16E : dout <= 12'hC41;
		12'h16F : dout <= 12'hC44;
		12'h170 : dout <= 12'hC47;
		12'h171 : dout <= 12'hC49;
		12'h172 : dout <= 12'hC4C;
		12'h173 : dout <= 12'hC4F;
		12'h174 : dout <= 12'hC51;
		12'h175 : dout <= 12'hC54;
		12'h176 : dout <= 12'hC57;
		12'h177 : dout <= 12'hC59;
		12'h178 : dout <= 12'hC5C;
		12'h179 : dout <= 12'hC5E;
		12'h17A : dout <= 12'hC61;
		12'h17B : dout <= 12'hC64;
		12'h17C : dout <= 12'hC66;
		12'h17D : dout <= 12'hC69;
		12'h17E : dout <= 12'hC6C;
		12'h17F : dout <= 12'hC6E;
		12'h180 : dout <= 12'hC71;
		12'h181 : dout <= 12'hC73;
		12'h182 : dout <= 12'hC76;
		12'h183 : dout <= 12'hC79;
		12'h184 : dout <= 12'hC7B;
		12'h185 : dout <= 12'hC7E;
		12'h186 : dout <= 12'hC80;
		12'h187 : dout <= 12'hC83;
		12'h188 : dout <= 12'hC86;
		12'h189 : dout <= 12'hC88;
		12'h18A : dout <= 12'hC8B;
		12'h18B : dout <= 12'hC8D;
		12'h18C : dout <= 12'hC90;
		12'h18D : dout <= 12'hC92;
		12'h18E : dout <= 12'hC95;
		12'h18F : dout <= 12'hC98;
		12'h190 : dout <= 12'hC9A;
		12'h191 : dout <= 12'hC9D;
		12'h192 : dout <= 12'hC9F;
		12'h193 : dout <= 12'hCA2;
		12'h194 : dout <= 12'hCA4;
		12'h195 : dout <= 12'hCA7;
		12'h196 : dout <= 12'hCAA;
		12'h197 : dout <= 12'hCAC;
		12'h198 : dout <= 12'hCAF;
		12'h199 : dout <= 12'hCB1;
		12'h19A : dout <= 12'hCB4;
		12'h19B : dout <= 12'hCB6;
		12'h19C : dout <= 12'hCB9;
		12'h19D : dout <= 12'hCBB;
		12'h19E : dout <= 12'hCBE;
		12'h19F : dout <= 12'hCC0;
		12'h1A0 : dout <= 12'hCC3;
		12'h1A1 : dout <= 12'hCC5;
		12'h1A2 : dout <= 12'hCC8;
		12'h1A3 : dout <= 12'hCCA;
		12'h1A4 : dout <= 12'hCCD;
		12'h1A5 : dout <= 12'hCCF;
		12'h1A6 : dout <= 12'hCD2;
		12'h1A7 : dout <= 12'hCD4;
		12'h1A8 : dout <= 12'hCD7;
		12'h1A9 : dout <= 12'hCD9;
		12'h1AA : dout <= 12'hCDC;
		12'h1AB : dout <= 12'hCDE;
		12'h1AC : dout <= 12'hCE1;
		12'h1AD : dout <= 12'hCE3;
		12'h1AE : dout <= 12'hCE6;
		12'h1AF : dout <= 12'hCE8;
		12'h1B0 : dout <= 12'hCEB;
		12'h1B1 : dout <= 12'hCED;
		12'h1B2 : dout <= 12'hCF0;
		12'h1B3 : dout <= 12'hCF2;
		12'h1B4 : dout <= 12'hCF5;
		12'h1B5 : dout <= 12'hCF7;
		12'h1B6 : dout <= 12'hCFA;
		12'h1B7 : dout <= 12'hCFC;
		12'h1B8 : dout <= 12'hCFF;
		12'h1B9 : dout <= 12'hD01;
		12'h1BA : dout <= 12'hD03;
		12'h1BB : dout <= 12'hD06;
		12'h1BC : dout <= 12'hD08;
		12'h1BD : dout <= 12'hD0B;
		12'h1BE : dout <= 12'hD0D;
		12'h1BF : dout <= 12'hD10;
		12'h1C0 : dout <= 12'hD12;
		12'h1C1 : dout <= 12'hD15;
		12'h1C2 : dout <= 12'hD17;
		12'h1C3 : dout <= 12'hD19;
		12'h1C4 : dout <= 12'hD1C;
		12'h1C5 : dout <= 12'hD1E;
		12'h1C6 : dout <= 12'hD21;
		12'h1C7 : dout <= 12'hD23;
		12'h1C8 : dout <= 12'hD25;
		12'h1C9 : dout <= 12'hD28;
		12'h1CA : dout <= 12'hD2A;
		12'h1CB : dout <= 12'hD2D;
		12'h1CC : dout <= 12'hD2F;
		12'h1CD : dout <= 12'hD31;
		12'h1CE : dout <= 12'hD34;
		12'h1CF : dout <= 12'hD36;
		12'h1D0 : dout <= 12'hD39;
		12'h1D1 : dout <= 12'hD3B;
		12'h1D2 : dout <= 12'hD3D;
		12'h1D3 : dout <= 12'hD40;
		12'h1D4 : dout <= 12'hD42;
		12'h1D5 : dout <= 12'hD44;
		12'h1D6 : dout <= 12'hD47;
		12'h1D7 : dout <= 12'hD49;
		12'h1D8 : dout <= 12'hD4B;
		12'h1D9 : dout <= 12'hD4E;
		12'h1DA : dout <= 12'hD50;
		12'h1DB : dout <= 12'hD53;
		12'h1DC : dout <= 12'hD55;
		12'h1DD : dout <= 12'hD57;
		12'h1DE : dout <= 12'hD5A;
		12'h1DF : dout <= 12'hD5C;
		12'h1E0 : dout <= 12'hD5E;
		12'h1E1 : dout <= 12'hD61;
		12'h1E2 : dout <= 12'hD63;
		12'h1E3 : dout <= 12'hD65;
		12'h1E4 : dout <= 12'hD67;
		12'h1E5 : dout <= 12'hD6A;
		12'h1E6 : dout <= 12'hD6C;
		12'h1E7 : dout <= 12'hD6E;
		12'h1E8 : dout <= 12'hD71;
		12'h1E9 : dout <= 12'hD73;
		12'h1EA : dout <= 12'hD75;
		12'h1EB : dout <= 12'hD78;
		12'h1EC : dout <= 12'hD7A;
		12'h1ED : dout <= 12'hD7C;
		12'h1EE : dout <= 12'hD7E;
		12'h1EF : dout <= 12'hD81;
		12'h1F0 : dout <= 12'hD83;
		12'h1F1 : dout <= 12'hD85;
		12'h1F2 : dout <= 12'hD88;
		12'h1F3 : dout <= 12'hD8A;
		12'h1F4 : dout <= 12'hD8C;
		12'h1F5 : dout <= 12'hD8E;
		12'h1F6 : dout <= 12'hD91;
		12'h1F7 : dout <= 12'hD93;
		12'h1F8 : dout <= 12'hD95;
		12'h1F9 : dout <= 12'hD97;
		12'h1FA : dout <= 12'hD9A;
		12'h1FB : dout <= 12'hD9C;
		12'h1FC : dout <= 12'hD9E;
		12'h1FD : dout <= 12'hDA0;
		12'h1FE : dout <= 12'hDA3;
		12'h1FF : dout <= 12'hDA5;
		12'h200 : dout <= 12'hDA7;
		12'h201 : dout <= 12'hDA9;
		12'h202 : dout <= 12'hDAB;
		12'h203 : dout <= 12'hDAE;
		12'h204 : dout <= 12'hDB0;
		12'h205 : dout <= 12'hDB2;
		12'h206 : dout <= 12'hDB4;
		12'h207 : dout <= 12'hDB6;
		12'h208 : dout <= 12'hDB9;
		12'h209 : dout <= 12'hDBB;
		12'h20A : dout <= 12'hDBD;
		12'h20B : dout <= 12'hDBF;
		12'h20C : dout <= 12'hDC1;
		12'h20D : dout <= 12'hDC4;
		12'h20E : dout <= 12'hDC6;
		12'h20F : dout <= 12'hDC8;
		12'h210 : dout <= 12'hDCA;
		12'h211 : dout <= 12'hDCC;
		12'h212 : dout <= 12'hDCE;
		12'h213 : dout <= 12'hDD1;
		12'h214 : dout <= 12'hDD3;
		12'h215 : dout <= 12'hDD5;
		12'h216 : dout <= 12'hDD7;
		12'h217 : dout <= 12'hDD9;
		12'h218 : dout <= 12'hDDB;
		12'h219 : dout <= 12'hDDD;
		12'h21A : dout <= 12'hDE0;
		12'h21B : dout <= 12'hDE2;
		12'h21C : dout <= 12'hDE4;
		12'h21D : dout <= 12'hDE6;
		12'h21E : dout <= 12'hDE8;
		12'h21F : dout <= 12'hDEA;
		12'h220 : dout <= 12'hDEC;
		12'h221 : dout <= 12'hDEE;
		12'h222 : dout <= 12'hDF0;
		12'h223 : dout <= 12'hDF3;
		12'h224 : dout <= 12'hDF5;
		12'h225 : dout <= 12'hDF7;
		12'h226 : dout <= 12'hDF9;
		12'h227 : dout <= 12'hDFB;
		12'h228 : dout <= 12'hDFD;
		12'h229 : dout <= 12'hDFF;
		12'h22A : dout <= 12'hE01;
		12'h22B : dout <= 12'hE03;
		12'h22C : dout <= 12'hE05;
		12'h22D : dout <= 12'hE07;
		12'h22E : dout <= 12'hE09;
		12'h22F : dout <= 12'hE0B;
		12'h230 : dout <= 12'hE0E;
		12'h231 : dout <= 12'hE10;
		12'h232 : dout <= 12'hE12;
		12'h233 : dout <= 12'hE14;
		12'h234 : dout <= 12'hE16;
		12'h235 : dout <= 12'hE18;
		12'h236 : dout <= 12'hE1A;
		12'h237 : dout <= 12'hE1C;
		12'h238 : dout <= 12'hE1E;
		12'h239 : dout <= 12'hE20;
		12'h23A : dout <= 12'hE22;
		12'h23B : dout <= 12'hE24;
		12'h23C : dout <= 12'hE26;
		12'h23D : dout <= 12'hE28;
		12'h23E : dout <= 12'hE2A;
		12'h23F : dout <= 12'hE2C;
		12'h240 : dout <= 12'hE2E;
		12'h241 : dout <= 12'hE30;
		12'h242 : dout <= 12'hE32;
		12'h243 : dout <= 12'hE34;
		12'h244 : dout <= 12'hE36;
		12'h245 : dout <= 12'hE38;
		12'h246 : dout <= 12'hE3A;
		12'h247 : dout <= 12'hE3C;
		12'h248 : dout <= 12'hE3E;
		12'h249 : dout <= 12'hE40;
		12'h24A : dout <= 12'hE42;
		12'h24B : dout <= 12'hE44;
		12'h24C : dout <= 12'hE45;
		12'h24D : dout <= 12'hE47;
		12'h24E : dout <= 12'hE49;
		12'h24F : dout <= 12'hE4B;
		12'h250 : dout <= 12'hE4D;
		12'h251 : dout <= 12'hE4F;
		12'h252 : dout <= 12'hE51;
		12'h253 : dout <= 12'hE53;
		12'h254 : dout <= 12'hE55;
		12'h255 : dout <= 12'hE57;
		12'h256 : dout <= 12'hE59;
		12'h257 : dout <= 12'hE5B;
		12'h258 : dout <= 12'hE5D;
		12'h259 : dout <= 12'hE5E;
		12'h25A : dout <= 12'hE60;
		12'h25B : dout <= 12'hE62;
		12'h25C : dout <= 12'hE64;
		12'h25D : dout <= 12'hE66;
		12'h25E : dout <= 12'hE68;
		12'h25F : dout <= 12'hE6A;
		12'h260 : dout <= 12'hE6C;
		12'h261 : dout <= 12'hE6E;
		12'h262 : dout <= 12'hE6F;
		12'h263 : dout <= 12'hE71;
		12'h264 : dout <= 12'hE73;
		12'h265 : dout <= 12'hE75;
		12'h266 : dout <= 12'hE77;
		12'h267 : dout <= 12'hE79;
		12'h268 : dout <= 12'hE7B;
		12'h269 : dout <= 12'hE7C;
		12'h26A : dout <= 12'hE7E;
		12'h26B : dout <= 12'hE80;
		12'h26C : dout <= 12'hE82;
		12'h26D : dout <= 12'hE84;
		12'h26E : dout <= 12'hE85;
		12'h26F : dout <= 12'hE87;
		12'h270 : dout <= 12'hE89;
		12'h271 : dout <= 12'hE8B;
		12'h272 : dout <= 12'hE8D;
		12'h273 : dout <= 12'hE8F;
		12'h274 : dout <= 12'hE90;
		12'h275 : dout <= 12'hE92;
		12'h276 : dout <= 12'hE94;
		12'h277 : dout <= 12'hE96;
		12'h278 : dout <= 12'hE97;
		12'h279 : dout <= 12'hE99;
		12'h27A : dout <= 12'hE9B;
		12'h27B : dout <= 12'hE9D;
		12'h27C : dout <= 12'hE9F;
		12'h27D : dout <= 12'hEA0;
		12'h27E : dout <= 12'hEA2;
		12'h27F : dout <= 12'hEA4;
		12'h280 : dout <= 12'hEA6;
		12'h281 : dout <= 12'hEA7;
		12'h282 : dout <= 12'hEA9;
		12'h283 : dout <= 12'hEAB;
		12'h284 : dout <= 12'hEAC;
		12'h285 : dout <= 12'hEAE;
		12'h286 : dout <= 12'hEB0;
		12'h287 : dout <= 12'hEB2;
		12'h288 : dout <= 12'hEB3;
		12'h289 : dout <= 12'hEB5;
		12'h28A : dout <= 12'hEB7;
		12'h28B : dout <= 12'hEB8;
		12'h28C : dout <= 12'hEBA;
		12'h28D : dout <= 12'hEBC;
		12'h28E : dout <= 12'hEBE;
		12'h28F : dout <= 12'hEBF;
		12'h290 : dout <= 12'hEC1;
		12'h291 : dout <= 12'hEC3;
		12'h292 : dout <= 12'hEC4;
		12'h293 : dout <= 12'hEC6;
		12'h294 : dout <= 12'hEC8;
		12'h295 : dout <= 12'hEC9;
		12'h296 : dout <= 12'hECB;
		12'h297 : dout <= 12'hECD;
		12'h298 : dout <= 12'hECE;
		12'h299 : dout <= 12'hED0;
		12'h29A : dout <= 12'hED2;
		12'h29B : dout <= 12'hED3;
		12'h29C : dout <= 12'hED5;
		12'h29D : dout <= 12'hED6;
		12'h29E : dout <= 12'hED8;
		12'h29F : dout <= 12'hEDA;
		12'h2A0 : dout <= 12'hEDB;
		12'h2A1 : dout <= 12'hEDD;
		12'h2A2 : dout <= 12'hEDE;
		12'h2A3 : dout <= 12'hEE0;
		12'h2A4 : dout <= 12'hEE2;
		12'h2A5 : dout <= 12'hEE3;
		12'h2A6 : dout <= 12'hEE5;
		12'h2A7 : dout <= 12'hEE6;
		12'h2A8 : dout <= 12'hEE8;
		12'h2A9 : dout <= 12'hEEA;
		12'h2AA : dout <= 12'hEEB;
		12'h2AB : dout <= 12'hEED;
		12'h2AC : dout <= 12'hEEE;
		12'h2AD : dout <= 12'hEF0;
		12'h2AE : dout <= 12'hEF1;
		12'h2AF : dout <= 12'hEF3;
		12'h2B0 : dout <= 12'hEF5;
		12'h2B1 : dout <= 12'hEF6;
		12'h2B2 : dout <= 12'hEF8;
		12'h2B3 : dout <= 12'hEF9;
		12'h2B4 : dout <= 12'hEFB;
		12'h2B5 : dout <= 12'hEFC;
		12'h2B6 : dout <= 12'hEFE;
		12'h2B7 : dout <= 12'hEFF;
		12'h2B8 : dout <= 12'hF01;
		12'h2B9 : dout <= 12'hF02;
		12'h2BA : dout <= 12'hF04;
		12'h2BB : dout <= 12'hF05;
		12'h2BC : dout <= 12'hF07;
		12'h2BD : dout <= 12'hF08;
		12'h2BE : dout <= 12'hF0A;
		12'h2BF : dout <= 12'hF0B;
		12'h2C0 : dout <= 12'hF0D;
		12'h2C1 : dout <= 12'hF0E;
		12'h2C2 : dout <= 12'hF10;
		12'h2C3 : dout <= 12'hF11;
		12'h2C4 : dout <= 12'hF13;
		12'h2C5 : dout <= 12'hF14;
		12'h2C6 : dout <= 12'hF16;
		12'h2C7 : dout <= 12'hF17;
		12'h2C8 : dout <= 12'hF18;
		12'h2C9 : dout <= 12'hF1A;
		12'h2CA : dout <= 12'hF1B;
		12'h2CB : dout <= 12'hF1D;
		12'h2CC : dout <= 12'hF1E;
		12'h2CD : dout <= 12'hF20;
		12'h2CE : dout <= 12'hF21;
		12'h2CF : dout <= 12'hF23;
		12'h2D0 : dout <= 12'hF24;
		12'h2D1 : dout <= 12'hF25;
		12'h2D2 : dout <= 12'hF27;
		12'h2D3 : dout <= 12'hF28;
		12'h2D4 : dout <= 12'hF2A;
		12'h2D5 : dout <= 12'hF2B;
		12'h2D6 : dout <= 12'hF2C;
		12'h2D7 : dout <= 12'hF2E;
		12'h2D8 : dout <= 12'hF2F;
		12'h2D9 : dout <= 12'hF30;
		12'h2DA : dout <= 12'hF32;
		12'h2DB : dout <= 12'hF33;
		12'h2DC : dout <= 12'hF35;
		12'h2DD : dout <= 12'hF36;
		12'h2DE : dout <= 12'hF37;
		12'h2DF : dout <= 12'hF39;
		12'h2E0 : dout <= 12'hF3A;
		12'h2E1 : dout <= 12'hF3B;
		12'h2E2 : dout <= 12'hF3D;
		12'h2E3 : dout <= 12'hF3E;
		12'h2E4 : dout <= 12'hF3F;
		12'h2E5 : dout <= 12'hF41;
		12'h2E6 : dout <= 12'hF42;
		12'h2E7 : dout <= 12'hF43;
		12'h2E8 : dout <= 12'hF45;
		12'h2E9 : dout <= 12'hF46;
		12'h2EA : dout <= 12'hF47;
		12'h2EB : dout <= 12'hF48;
		12'h2EC : dout <= 12'hF4A;
		12'h2ED : dout <= 12'hF4B;
		12'h2EE : dout <= 12'hF4C;
		12'h2EF : dout <= 12'hF4E;
		12'h2F0 : dout <= 12'hF4F;
		12'h2F1 : dout <= 12'hF50;
		12'h2F2 : dout <= 12'hF51;
		12'h2F3 : dout <= 12'hF53;
		12'h2F4 : dout <= 12'hF54;
		12'h2F5 : dout <= 12'hF55;
		12'h2F6 : dout <= 12'hF56;
		12'h2F7 : dout <= 12'hF58;
		12'h2F8 : dout <= 12'hF59;
		12'h2F9 : dout <= 12'hF5A;
		12'h2FA : dout <= 12'hF5B;
		12'h2FB : dout <= 12'hF5D;
		12'h2FC : dout <= 12'hF5E;
		12'h2FD : dout <= 12'hF5F;
		12'h2FE : dout <= 12'hF60;
		12'h2FF : dout <= 12'hF61;
		12'h300 : dout <= 12'hF63;
		12'h301 : dout <= 12'hF64;
		12'h302 : dout <= 12'hF65;
		12'h303 : dout <= 12'hF66;
		12'h304 : dout <= 12'hF67;
		12'h305 : dout <= 12'hF69;
		12'h306 : dout <= 12'hF6A;
		12'h307 : dout <= 12'hF6B;
		12'h308 : dout <= 12'hF6C;
		12'h309 : dout <= 12'hF6D;
		12'h30A : dout <= 12'hF6E;
		12'h30B : dout <= 12'hF70;
		12'h30C : dout <= 12'hF71;
		12'h30D : dout <= 12'hF72;
		12'h30E : dout <= 12'hF73;
		12'h30F : dout <= 12'hF74;
		12'h310 : dout <= 12'hF75;
		12'h311 : dout <= 12'hF76;
		12'h312 : dout <= 12'hF78;
		12'h313 : dout <= 12'hF79;
		12'h314 : dout <= 12'hF7A;
		12'h315 : dout <= 12'hF7B;
		12'h316 : dout <= 12'hF7C;
		12'h317 : dout <= 12'hF7D;
		12'h318 : dout <= 12'hF7E;
		12'h319 : dout <= 12'hF7F;
		12'h31A : dout <= 12'hF80;
		12'h31B : dout <= 12'hF81;
		12'h31C : dout <= 12'hF83;
		12'h31D : dout <= 12'hF84;
		12'h31E : dout <= 12'hF85;
		12'h31F : dout <= 12'hF86;
		12'h320 : dout <= 12'hF87;
		12'h321 : dout <= 12'hF88;
		12'h322 : dout <= 12'hF89;
		12'h323 : dout <= 12'hF8A;
		12'h324 : dout <= 12'hF8B;
		12'h325 : dout <= 12'hF8C;
		12'h326 : dout <= 12'hF8D;
		12'h327 : dout <= 12'hF8E;
		12'h328 : dout <= 12'hF8F;
		12'h329 : dout <= 12'hF90;
		12'h32A : dout <= 12'hF91;
		12'h32B : dout <= 12'hF92;
		12'h32C : dout <= 12'hF93;
		12'h32D : dout <= 12'hF94;
		12'h32E : dout <= 12'hF95;
		12'h32F : dout <= 12'hF96;
		12'h330 : dout <= 12'hF97;
		12'h331 : dout <= 12'hF98;
		12'h332 : dout <= 12'hF99;
		12'h333 : dout <= 12'hF9A;
		12'h334 : dout <= 12'hF9B;
		12'h335 : dout <= 12'hF9C;
		12'h336 : dout <= 12'hF9D;
		12'h337 : dout <= 12'hF9E;
		12'h338 : dout <= 12'hF9F;
		12'h339 : dout <= 12'hFA0;
		12'h33A : dout <= 12'hFA1;
		12'h33B : dout <= 12'hFA2;
		12'h33C : dout <= 12'hFA3;
		12'h33D : dout <= 12'hFA4;
		12'h33E : dout <= 12'hFA5;
		12'h33F : dout <= 12'hFA5;
		12'h340 : dout <= 12'hFA6;
		12'h341 : dout <= 12'hFA7;
		12'h342 : dout <= 12'hFA8;
		12'h343 : dout <= 12'hFA9;
		12'h344 : dout <= 12'hFAA;
		12'h345 : dout <= 12'hFAB;
		12'h346 : dout <= 12'hFAC;
		12'h347 : dout <= 12'hFAD;
		12'h348 : dout <= 12'hFAE;
		12'h349 : dout <= 12'hFAE;
		12'h34A : dout <= 12'hFAF;
		12'h34B : dout <= 12'hFB0;
		12'h34C : dout <= 12'hFB1;
		12'h34D : dout <= 12'hFB2;
		12'h34E : dout <= 12'hFB3;
		12'h34F : dout <= 12'hFB4;
		12'h350 : dout <= 12'hFB4;
		12'h351 : dout <= 12'hFB5;
		12'h352 : dout <= 12'hFB6;
		12'h353 : dout <= 12'hFB7;
		12'h354 : dout <= 12'hFB8;
		12'h355 : dout <= 12'hFB8;
		12'h356 : dout <= 12'hFB9;
		12'h357 : dout <= 12'hFBA;
		12'h358 : dout <= 12'hFBB;
		12'h359 : dout <= 12'hFBC;
		12'h35A : dout <= 12'hFBC;
		12'h35B : dout <= 12'hFBD;
		12'h35C : dout <= 12'hFBE;
		12'h35D : dout <= 12'hFBF;
		12'h35E : dout <= 12'hFC0;
		12'h35F : dout <= 12'hFC0;
		12'h360 : dout <= 12'hFC1;
		12'h361 : dout <= 12'hFC2;
		12'h362 : dout <= 12'hFC3;
		12'h363 : dout <= 12'hFC3;
		12'h364 : dout <= 12'hFC4;
		12'h365 : dout <= 12'hFC5;
		12'h366 : dout <= 12'hFC6;
		12'h367 : dout <= 12'hFC6;
		12'h368 : dout <= 12'hFC7;
		12'h369 : dout <= 12'hFC8;
		12'h36A : dout <= 12'hFC9;
		12'h36B : dout <= 12'hFC9;
		12'h36C : dout <= 12'hFCA;
		12'h36D : dout <= 12'hFCB;
		12'h36E : dout <= 12'hFCB;
		12'h36F : dout <= 12'hFCC;
		12'h370 : dout <= 12'hFCD;
		12'h371 : dout <= 12'hFCD;
		12'h372 : dout <= 12'hFCE;
		12'h373 : dout <= 12'hFCF;
		12'h374 : dout <= 12'hFCF;
		12'h375 : dout <= 12'hFD0;
		12'h376 : dout <= 12'hFD1;
		12'h377 : dout <= 12'hFD1;
		12'h378 : dout <= 12'hFD2;
		12'h379 : dout <= 12'hFD3;
		12'h37A : dout <= 12'hFD3;
		12'h37B : dout <= 12'hFD4;
		12'h37C : dout <= 12'hFD5;
		12'h37D : dout <= 12'hFD5;
		12'h37E : dout <= 12'hFD6;
		12'h37F : dout <= 12'hFD7;
		12'h380 : dout <= 12'hFD7;
		12'h381 : dout <= 12'hFD8;
		12'h382 : dout <= 12'hFD8;
		12'h383 : dout <= 12'hFD9;
		12'h384 : dout <= 12'hFDA;
		12'h385 : dout <= 12'hFDA;
		12'h386 : dout <= 12'hFDB;
		12'h387 : dout <= 12'hFDB;
		12'h388 : dout <= 12'hFDC;
		12'h389 : dout <= 12'hFDC;
		12'h38A : dout <= 12'hFDD;
		12'h38B : dout <= 12'hFDE;
		12'h38C : dout <= 12'hFDE;
		12'h38D : dout <= 12'hFDF;
		12'h38E : dout <= 12'hFDF;
		12'h38F : dout <= 12'hFE0;
		12'h390 : dout <= 12'hFE0;
		12'h391 : dout <= 12'hFE1;
		12'h392 : dout <= 12'hFE1;
		12'h393 : dout <= 12'hFE2;
		12'h394 : dout <= 12'hFE2;
		12'h395 : dout <= 12'hFE3;
		12'h396 : dout <= 12'hFE3;
		12'h397 : dout <= 12'hFE4;
		12'h398 : dout <= 12'hFE5;
		12'h399 : dout <= 12'hFE5;
		12'h39A : dout <= 12'hFE5;
		12'h39B : dout <= 12'hFE6;
		12'h39C : dout <= 12'hFE6;
		12'h39D : dout <= 12'hFE7;
		12'h39E : dout <= 12'hFE7;
		12'h39F : dout <= 12'hFE8;
		12'h3A0 : dout <= 12'hFE8;
		12'h3A1 : dout <= 12'hFE9;
		12'h3A2 : dout <= 12'hFE9;
		12'h3A3 : dout <= 12'hFEA;
		12'h3A4 : dout <= 12'hFEA;
		12'h3A5 : dout <= 12'hFEB;
		12'h3A6 : dout <= 12'hFEB;
		12'h3A7 : dout <= 12'hFEB;
		12'h3A8 : dout <= 12'hFEC;
		12'h3A9 : dout <= 12'hFEC;
		12'h3AA : dout <= 12'hFED;
		12'h3AB : dout <= 12'hFED;
		12'h3AC : dout <= 12'hFEE;
		12'h3AD : dout <= 12'hFEE;
		12'h3AE : dout <= 12'hFEE;
		12'h3AF : dout <= 12'hFEF;
		12'h3B0 : dout <= 12'hFEF;
		12'h3B1 : dout <= 12'hFEF;
		12'h3B2 : dout <= 12'hFF0;
		12'h3B3 : dout <= 12'hFF0;
		12'h3B4 : dout <= 12'hFF1;
		12'h3B5 : dout <= 12'hFF1;
		12'h3B6 : dout <= 12'hFF1;
		12'h3B7 : dout <= 12'hFF2;
		12'h3B8 : dout <= 12'hFF2;
		12'h3B9 : dout <= 12'hFF2;
		12'h3BA : dout <= 12'hFF3;
		12'h3BB : dout <= 12'hFF3;
		12'h3BC : dout <= 12'hFF3;
		12'h3BD : dout <= 12'hFF4;
		12'h3BE : dout <= 12'hFF4;
		12'h3BF : dout <= 12'hFF4;
		12'h3C0 : dout <= 12'hFF5;
		12'h3C1 : dout <= 12'hFF5;
		12'h3C2 : dout <= 12'hFF5;
		12'h3C3 : dout <= 12'hFF6;
		12'h3C4 : dout <= 12'hFF6;
		12'h3C5 : dout <= 12'hFF6;
		12'h3C6 : dout <= 12'hFF6;
		12'h3C7 : dout <= 12'hFF7;
		12'h3C8 : dout <= 12'hFF7;
		12'h3C9 : dout <= 12'hFF7;
		12'h3CA : dout <= 12'hFF7;
		12'h3CB : dout <= 12'hFF8;
		12'h3CC : dout <= 12'hFF8;
		12'h3CD : dout <= 12'hFF8;
		12'h3CE : dout <= 12'hFF8;
		12'h3CF : dout <= 12'hFF9;
		12'h3D0 : dout <= 12'hFF9;
		12'h3D1 : dout <= 12'hFF9;
		12'h3D2 : dout <= 12'hFF9;
		12'h3D3 : dout <= 12'hFFA;
		12'h3D4 : dout <= 12'hFFA;
		12'h3D5 : dout <= 12'hFFA;
		12'h3D6 : dout <= 12'hFFA;
		12'h3D7 : dout <= 12'hFFA;
		12'h3D8 : dout <= 12'hFFB;
		12'h3D9 : dout <= 12'hFFB;
		12'h3DA : dout <= 12'hFFB;
		12'h3DB : dout <= 12'hFFB;
		12'h3DC : dout <= 12'hFFB;
		12'h3DD : dout <= 12'hFFC;
		12'h3DE : dout <= 12'hFFC;
		12'h3DF : dout <= 12'hFFC;
		12'h3E0 : dout <= 12'hFFC;
		12'h3E1 : dout <= 12'hFFC;
		12'h3E2 : dout <= 12'hFFC;
		12'h3E3 : dout <= 12'hFFC;
		12'h3E4 : dout <= 12'hFFD;
		12'h3E5 : dout <= 12'hFFD;
		12'h3E6 : dout <= 12'hFFD;
		12'h3E7 : dout <= 12'hFFD;
		12'h3E8 : dout <= 12'hFFD;
		12'h3E9 : dout <= 12'hFFD;
		12'h3EA : dout <= 12'hFFD;
		12'h3EB : dout <= 12'hFFD;
		12'h3EC : dout <= 12'hFFE;
		12'h3ED : dout <= 12'hFFE;
		12'h3EE : dout <= 12'hFFE;
		12'h3EF : dout <= 12'hFFE;
		12'h3F0 : dout <= 12'hFFE;
		12'h3F1 : dout <= 12'hFFE;
		12'h3F2 : dout <= 12'hFFE;
		12'h3F3 : dout <= 12'hFFE;
		12'h3F4 : dout <= 12'hFFE;
		12'h3F5 : dout <= 12'hFFE;
		12'h3F6 : dout <= 12'hFFE;
		12'h3F7 : dout <= 12'hFFE;
		12'h3F8 : dout <= 12'hFFE;
		12'h3F9 : dout <= 12'hFFE;
		12'h3FA : dout <= 12'hFFE;
		12'h3FB : dout <= 12'hFFE;
		12'h3FC : dout <= 12'hFFE;
		12'h3FD : dout <= 12'hFFE;
		12'h3FE : dout <= 12'hFFE;
		12'h3FF : dout <= 12'hFFE;
		12'h400 : dout <= 12'hFFF;
		12'h401 : dout <= 12'hFFE;
		12'h402 : dout <= 12'hFFE;
		12'h403 : dout <= 12'hFFE;
		12'h404 : dout <= 12'hFFE;
		12'h405 : dout <= 12'hFFE;
		12'h406 : dout <= 12'hFFE;
		12'h407 : dout <= 12'hFFE;
		12'h408 : dout <= 12'hFFE;
		12'h409 : dout <= 12'hFFE;
		12'h40A : dout <= 12'hFFE;
		12'h40B : dout <= 12'hFFE;
		12'h40C : dout <= 12'hFFE;
		12'h40D : dout <= 12'hFFE;
		12'h40E : dout <= 12'hFFE;
		12'h40F : dout <= 12'hFFE;
		12'h410 : dout <= 12'hFFE;
		12'h411 : dout <= 12'hFFE;
		12'h412 : dout <= 12'hFFE;
		12'h413 : dout <= 12'hFFE;
		12'h414 : dout <= 12'hFFE;
		12'h415 : dout <= 12'hFFD;
		12'h416 : dout <= 12'hFFD;
		12'h417 : dout <= 12'hFFD;
		12'h418 : dout <= 12'hFFD;
		12'h419 : dout <= 12'hFFD;
		12'h41A : dout <= 12'hFFD;
		12'h41B : dout <= 12'hFFD;
		12'h41C : dout <= 12'hFFD;
		12'h41D : dout <= 12'hFFC;
		12'h41E : dout <= 12'hFFC;
		12'h41F : dout <= 12'hFFC;
		12'h420 : dout <= 12'hFFC;
		12'h421 : dout <= 12'hFFC;
		12'h422 : dout <= 12'hFFC;
		12'h423 : dout <= 12'hFFC;
		12'h424 : dout <= 12'hFFB;
		12'h425 : dout <= 12'hFFB;
		12'h426 : dout <= 12'hFFB;
		12'h427 : dout <= 12'hFFB;
		12'h428 : dout <= 12'hFFB;
		12'h429 : dout <= 12'hFFA;
		12'h42A : dout <= 12'hFFA;
		12'h42B : dout <= 12'hFFA;
		12'h42C : dout <= 12'hFFA;
		12'h42D : dout <= 12'hFFA;
		12'h42E : dout <= 12'hFF9;
		12'h42F : dout <= 12'hFF9;
		12'h430 : dout <= 12'hFF9;
		12'h431 : dout <= 12'hFF9;
		12'h432 : dout <= 12'hFF8;
		12'h433 : dout <= 12'hFF8;
		12'h434 : dout <= 12'hFF8;
		12'h435 : dout <= 12'hFF8;
		12'h436 : dout <= 12'hFF7;
		12'h437 : dout <= 12'hFF7;
		12'h438 : dout <= 12'hFF7;
		12'h439 : dout <= 12'hFF7;
		12'h43A : dout <= 12'hFF6;
		12'h43B : dout <= 12'hFF6;
		12'h43C : dout <= 12'hFF6;
		12'h43D : dout <= 12'hFF6;
		12'h43E : dout <= 12'hFF5;
		12'h43F : dout <= 12'hFF5;
		12'h440 : dout <= 12'hFF5;
		12'h441 : dout <= 12'hFF4;
		12'h442 : dout <= 12'hFF4;
		12'h443 : dout <= 12'hFF4;
		12'h444 : dout <= 12'hFF3;
		12'h445 : dout <= 12'hFF3;
		12'h446 : dout <= 12'hFF3;
		12'h447 : dout <= 12'hFF2;
		12'h448 : dout <= 12'hFF2;
		12'h449 : dout <= 12'hFF2;
		12'h44A : dout <= 12'hFF1;
		12'h44B : dout <= 12'hFF1;
		12'h44C : dout <= 12'hFF1;
		12'h44D : dout <= 12'hFF0;
		12'h44E : dout <= 12'hFF0;
		12'h44F : dout <= 12'hFEF;
		12'h450 : dout <= 12'hFEF;
		12'h451 : dout <= 12'hFEF;
		12'h452 : dout <= 12'hFEE;
		12'h453 : dout <= 12'hFEE;
		12'h454 : dout <= 12'hFEE;
		12'h455 : dout <= 12'hFED;
		12'h456 : dout <= 12'hFED;
		12'h457 : dout <= 12'hFEC;
		12'h458 : dout <= 12'hFEC;
		12'h459 : dout <= 12'hFEB;
		12'h45A : dout <= 12'hFEB;
		12'h45B : dout <= 12'hFEB;
		12'h45C : dout <= 12'hFEA;
		12'h45D : dout <= 12'hFEA;
		12'h45E : dout <= 12'hFE9;
		12'h45F : dout <= 12'hFE9;
		12'h460 : dout <= 12'hFE8;
		12'h461 : dout <= 12'hFE8;
		12'h462 : dout <= 12'hFE7;
		12'h463 : dout <= 12'hFE7;
		12'h464 : dout <= 12'hFE6;
		12'h465 : dout <= 12'hFE6;
		12'h466 : dout <= 12'hFE5;
		12'h467 : dout <= 12'hFE5;
		12'h468 : dout <= 12'hFE5;
		12'h469 : dout <= 12'hFE4;
		12'h46A : dout <= 12'hFE3;
		12'h46B : dout <= 12'hFE3;
		12'h46C : dout <= 12'hFE2;
		12'h46D : dout <= 12'hFE2;
		12'h46E : dout <= 12'hFE1;
		12'h46F : dout <= 12'hFE1;
		12'h470 : dout <= 12'hFE0;
		12'h471 : dout <= 12'hFE0;
		12'h472 : dout <= 12'hFDF;
		12'h473 : dout <= 12'hFDF;
		12'h474 : dout <= 12'hFDE;
		12'h475 : dout <= 12'hFDE;
		12'h476 : dout <= 12'hFDD;
		12'h477 : dout <= 12'hFDC;
		12'h478 : dout <= 12'hFDC;
		12'h479 : dout <= 12'hFDB;
		12'h47A : dout <= 12'hFDB;
		12'h47B : dout <= 12'hFDA;
		12'h47C : dout <= 12'hFDA;
		12'h47D : dout <= 12'hFD9;
		12'h47E : dout <= 12'hFD8;
		12'h47F : dout <= 12'hFD8;
		12'h480 : dout <= 12'hFD7;
		12'h481 : dout <= 12'hFD7;
		12'h482 : dout <= 12'hFD6;
		12'h483 : dout <= 12'hFD5;
		12'h484 : dout <= 12'hFD5;
		12'h485 : dout <= 12'hFD4;
		12'h486 : dout <= 12'hFD3;
		12'h487 : dout <= 12'hFD3;
		12'h488 : dout <= 12'hFD2;
		12'h489 : dout <= 12'hFD1;
		12'h48A : dout <= 12'hFD1;
		12'h48B : dout <= 12'hFD0;
		12'h48C : dout <= 12'hFCF;
		12'h48D : dout <= 12'hFCF;
		12'h48E : dout <= 12'hFCE;
		12'h48F : dout <= 12'hFCD;
		12'h490 : dout <= 12'hFCD;
		12'h491 : dout <= 12'hFCC;
		12'h492 : dout <= 12'hFCB;
		12'h493 : dout <= 12'hFCB;
		12'h494 : dout <= 12'hFCA;
		12'h495 : dout <= 12'hFC9;
		12'h496 : dout <= 12'hFC9;
		12'h497 : dout <= 12'hFC8;
		12'h498 : dout <= 12'hFC7;
		12'h499 : dout <= 12'hFC6;
		12'h49A : dout <= 12'hFC6;
		12'h49B : dout <= 12'hFC5;
		12'h49C : dout <= 12'hFC4;
		12'h49D : dout <= 12'hFC3;
		12'h49E : dout <= 12'hFC3;
		12'h49F : dout <= 12'hFC2;
		12'h4A0 : dout <= 12'hFC1;
		12'h4A1 : dout <= 12'hFC0;
		12'h4A2 : dout <= 12'hFC0;
		12'h4A3 : dout <= 12'hFBF;
		12'h4A4 : dout <= 12'hFBE;
		12'h4A5 : dout <= 12'hFBD;
		12'h4A6 : dout <= 12'hFBC;
		12'h4A7 : dout <= 12'hFBC;
		12'h4A8 : dout <= 12'hFBB;
		12'h4A9 : dout <= 12'hFBA;
		12'h4AA : dout <= 12'hFB9;
		12'h4AB : dout <= 12'hFB8;
		12'h4AC : dout <= 12'hFB8;
		12'h4AD : dout <= 12'hFB7;
		12'h4AE : dout <= 12'hFB6;
		12'h4AF : dout <= 12'hFB5;
		12'h4B0 : dout <= 12'hFB4;
		12'h4B1 : dout <= 12'hFB4;
		12'h4B2 : dout <= 12'hFB3;
		12'h4B3 : dout <= 12'hFB2;
		12'h4B4 : dout <= 12'hFB1;
		12'h4B5 : dout <= 12'hFB0;
		12'h4B6 : dout <= 12'hFAF;
		12'h4B7 : dout <= 12'hFAE;
		12'h4B8 : dout <= 12'hFAE;
		12'h4B9 : dout <= 12'hFAD;
		12'h4BA : dout <= 12'hFAC;
		12'h4BB : dout <= 12'hFAB;
		12'h4BC : dout <= 12'hFAA;
		12'h4BD : dout <= 12'hFA9;
		12'h4BE : dout <= 12'hFA8;
		12'h4BF : dout <= 12'hFA7;
		12'h4C0 : dout <= 12'hFA6;
		12'h4C1 : dout <= 12'hFA5;
		12'h4C2 : dout <= 12'hFA5;
		12'h4C3 : dout <= 12'hFA4;
		12'h4C4 : dout <= 12'hFA3;
		12'h4C5 : dout <= 12'hFA2;
		12'h4C6 : dout <= 12'hFA1;
		12'h4C7 : dout <= 12'hFA0;
		12'h4C8 : dout <= 12'hF9F;
		12'h4C9 : dout <= 12'hF9E;
		12'h4CA : dout <= 12'hF9D;
		12'h4CB : dout <= 12'hF9C;
		12'h4CC : dout <= 12'hF9B;
		12'h4CD : dout <= 12'hF9A;
		12'h4CE : dout <= 12'hF99;
		12'h4CF : dout <= 12'hF98;
		12'h4D0 : dout <= 12'hF97;
		12'h4D1 : dout <= 12'hF96;
		12'h4D2 : dout <= 12'hF95;
		12'h4D3 : dout <= 12'hF94;
		12'h4D4 : dout <= 12'hF93;
		12'h4D5 : dout <= 12'hF92;
		12'h4D6 : dout <= 12'hF91;
		12'h4D7 : dout <= 12'hF90;
		12'h4D8 : dout <= 12'hF8F;
		12'h4D9 : dout <= 12'hF8E;
		12'h4DA : dout <= 12'hF8D;
		12'h4DB : dout <= 12'hF8C;
		12'h4DC : dout <= 12'hF8B;
		12'h4DD : dout <= 12'hF8A;
		12'h4DE : dout <= 12'hF89;
		12'h4DF : dout <= 12'hF88;
		12'h4E0 : dout <= 12'hF87;
		12'h4E1 : dout <= 12'hF86;
		12'h4E2 : dout <= 12'hF85;
		12'h4E3 : dout <= 12'hF84;
		12'h4E4 : dout <= 12'hF83;
		12'h4E5 : dout <= 12'hF81;
		12'h4E6 : dout <= 12'hF80;
		12'h4E7 : dout <= 12'hF7F;
		12'h4E8 : dout <= 12'hF7E;
		12'h4E9 : dout <= 12'hF7D;
		12'h4EA : dout <= 12'hF7C;
		12'h4EB : dout <= 12'hF7B;
		12'h4EC : dout <= 12'hF7A;
		12'h4ED : dout <= 12'hF79;
		12'h4EE : dout <= 12'hF78;
		12'h4EF : dout <= 12'hF76;
		12'h4F0 : dout <= 12'hF75;
		12'h4F1 : dout <= 12'hF74;
		12'h4F2 : dout <= 12'hF73;
		12'h4F3 : dout <= 12'hF72;
		12'h4F4 : dout <= 12'hF71;
		12'h4F5 : dout <= 12'hF70;
		12'h4F6 : dout <= 12'hF6E;
		12'h4F7 : dout <= 12'hF6D;
		12'h4F8 : dout <= 12'hF6C;
		12'h4F9 : dout <= 12'hF6B;
		12'h4FA : dout <= 12'hF6A;
		12'h4FB : dout <= 12'hF69;
		12'h4FC : dout <= 12'hF67;
		12'h4FD : dout <= 12'hF66;
		12'h4FE : dout <= 12'hF65;
		12'h4FF : dout <= 12'hF64;
		12'h500 : dout <= 12'hF63;
		12'h501 : dout <= 12'hF61;
		12'h502 : dout <= 12'hF60;
		12'h503 : dout <= 12'hF5F;
		12'h504 : dout <= 12'hF5E;
		12'h505 : dout <= 12'hF5D;
		12'h506 : dout <= 12'hF5B;
		12'h507 : dout <= 12'hF5A;
		12'h508 : dout <= 12'hF59;
		12'h509 : dout <= 12'hF58;
		12'h50A : dout <= 12'hF56;
		12'h50B : dout <= 12'hF55;
		12'h50C : dout <= 12'hF54;
		12'h50D : dout <= 12'hF53;
		12'h50E : dout <= 12'hF51;
		12'h50F : dout <= 12'hF50;
		12'h510 : dout <= 12'hF4F;
		12'h511 : dout <= 12'hF4E;
		12'h512 : dout <= 12'hF4C;
		12'h513 : dout <= 12'hF4B;
		12'h514 : dout <= 12'hF4A;
		12'h515 : dout <= 12'hF48;
		12'h516 : dout <= 12'hF47;
		12'h517 : dout <= 12'hF46;
		12'h518 : dout <= 12'hF45;
		12'h519 : dout <= 12'hF43;
		12'h51A : dout <= 12'hF42;
		12'h51B : dout <= 12'hF41;
		12'h51C : dout <= 12'hF3F;
		12'h51D : dout <= 12'hF3E;
		12'h51E : dout <= 12'hF3D;
		12'h51F : dout <= 12'hF3B;
		12'h520 : dout <= 12'hF3A;
		12'h521 : dout <= 12'hF39;
		12'h522 : dout <= 12'hF37;
		12'h523 : dout <= 12'hF36;
		12'h524 : dout <= 12'hF35;
		12'h525 : dout <= 12'hF33;
		12'h526 : dout <= 12'hF32;
		12'h527 : dout <= 12'hF30;
		12'h528 : dout <= 12'hF2F;
		12'h529 : dout <= 12'hF2E;
		12'h52A : dout <= 12'hF2C;
		12'h52B : dout <= 12'hF2B;
		12'h52C : dout <= 12'hF2A;
		12'h52D : dout <= 12'hF28;
		12'h52E : dout <= 12'hF27;
		12'h52F : dout <= 12'hF25;
		12'h530 : dout <= 12'hF24;
		12'h531 : dout <= 12'hF23;
		12'h532 : dout <= 12'hF21;
		12'h533 : dout <= 12'hF20;
		12'h534 : dout <= 12'hF1E;
		12'h535 : dout <= 12'hF1D;
		12'h536 : dout <= 12'hF1B;
		12'h537 : dout <= 12'hF1A;
		12'h538 : dout <= 12'hF18;
		12'h539 : dout <= 12'hF17;
		12'h53A : dout <= 12'hF16;
		12'h53B : dout <= 12'hF14;
		12'h53C : dout <= 12'hF13;
		12'h53D : dout <= 12'hF11;
		12'h53E : dout <= 12'hF10;
		12'h53F : dout <= 12'hF0E;
		12'h540 : dout <= 12'hF0D;
		12'h541 : dout <= 12'hF0B;
		12'h542 : dout <= 12'hF0A;
		12'h543 : dout <= 12'hF08;
		12'h544 : dout <= 12'hF07;
		12'h545 : dout <= 12'hF05;
		12'h546 : dout <= 12'hF04;
		12'h547 : dout <= 12'hF02;
		12'h548 : dout <= 12'hF01;
		12'h549 : dout <= 12'hEFF;
		12'h54A : dout <= 12'hEFE;
		12'h54B : dout <= 12'hEFC;
		12'h54C : dout <= 12'hEFB;
		12'h54D : dout <= 12'hEF9;
		12'h54E : dout <= 12'hEF8;
		12'h54F : dout <= 12'hEF6;
		12'h550 : dout <= 12'hEF5;
		12'h551 : dout <= 12'hEF3;
		12'h552 : dout <= 12'hEF1;
		12'h553 : dout <= 12'hEF0;
		12'h554 : dout <= 12'hEEE;
		12'h555 : dout <= 12'hEED;
		12'h556 : dout <= 12'hEEB;
		12'h557 : dout <= 12'hEEA;
		12'h558 : dout <= 12'hEE8;
		12'h559 : dout <= 12'hEE6;
		12'h55A : dout <= 12'hEE5;
		12'h55B : dout <= 12'hEE3;
		12'h55C : dout <= 12'hEE2;
		12'h55D : dout <= 12'hEE0;
		12'h55E : dout <= 12'hEDE;
		12'h55F : dout <= 12'hEDD;
		12'h560 : dout <= 12'hEDB;
		12'h561 : dout <= 12'hEDA;
		12'h562 : dout <= 12'hED8;
		12'h563 : dout <= 12'hED6;
		12'h564 : dout <= 12'hED5;
		12'h565 : dout <= 12'hED3;
		12'h566 : dout <= 12'hED2;
		12'h567 : dout <= 12'hED0;
		12'h568 : dout <= 12'hECE;
		12'h569 : dout <= 12'hECD;
		12'h56A : dout <= 12'hECB;
		12'h56B : dout <= 12'hEC9;
		12'h56C : dout <= 12'hEC8;
		12'h56D : dout <= 12'hEC6;
		12'h56E : dout <= 12'hEC4;
		12'h56F : dout <= 12'hEC3;
		12'h570 : dout <= 12'hEC1;
		12'h571 : dout <= 12'hEBF;
		12'h572 : dout <= 12'hEBE;
		12'h573 : dout <= 12'hEBC;
		12'h574 : dout <= 12'hEBA;
		12'h575 : dout <= 12'hEB8;
		12'h576 : dout <= 12'hEB7;
		12'h577 : dout <= 12'hEB5;
		12'h578 : dout <= 12'hEB3;
		12'h579 : dout <= 12'hEB2;
		12'h57A : dout <= 12'hEB0;
		12'h57B : dout <= 12'hEAE;
		12'h57C : dout <= 12'hEAC;
		12'h57D : dout <= 12'hEAB;
		12'h57E : dout <= 12'hEA9;
		12'h57F : dout <= 12'hEA7;
		12'h580 : dout <= 12'hEA6;
		12'h581 : dout <= 12'hEA4;
		12'h582 : dout <= 12'hEA2;
		12'h583 : dout <= 12'hEA0;
		12'h584 : dout <= 12'hE9F;
		12'h585 : dout <= 12'hE9D;
		12'h586 : dout <= 12'hE9B;
		12'h587 : dout <= 12'hE99;
		12'h588 : dout <= 12'hE97;
		12'h589 : dout <= 12'hE96;
		12'h58A : dout <= 12'hE94;
		12'h58B : dout <= 12'hE92;
		12'h58C : dout <= 12'hE90;
		12'h58D : dout <= 12'hE8F;
		12'h58E : dout <= 12'hE8D;
		12'h58F : dout <= 12'hE8B;
		12'h590 : dout <= 12'hE89;
		12'h591 : dout <= 12'hE87;
		12'h592 : dout <= 12'hE85;
		12'h593 : dout <= 12'hE84;
		12'h594 : dout <= 12'hE82;
		12'h595 : dout <= 12'hE80;
		12'h596 : dout <= 12'hE7E;
		12'h597 : dout <= 12'hE7C;
		12'h598 : dout <= 12'hE7B;
		12'h599 : dout <= 12'hE79;
		12'h59A : dout <= 12'hE77;
		12'h59B : dout <= 12'hE75;
		12'h59C : dout <= 12'hE73;
		12'h59D : dout <= 12'hE71;
		12'h59E : dout <= 12'hE6F;
		12'h59F : dout <= 12'hE6E;
		12'h5A0 : dout <= 12'hE6C;
		12'h5A1 : dout <= 12'hE6A;
		12'h5A2 : dout <= 12'hE68;
		12'h5A3 : dout <= 12'hE66;
		12'h5A4 : dout <= 12'hE64;
		12'h5A5 : dout <= 12'hE62;
		12'h5A6 : dout <= 12'hE60;
		12'h5A7 : dout <= 12'hE5E;
		12'h5A8 : dout <= 12'hE5D;
		12'h5A9 : dout <= 12'hE5B;
		12'h5AA : dout <= 12'hE59;
		12'h5AB : dout <= 12'hE57;
		12'h5AC : dout <= 12'hE55;
		12'h5AD : dout <= 12'hE53;
		12'h5AE : dout <= 12'hE51;
		12'h5AF : dout <= 12'hE4F;
		12'h5B0 : dout <= 12'hE4D;
		12'h5B1 : dout <= 12'hE4B;
		12'h5B2 : dout <= 12'hE49;
		12'h5B3 : dout <= 12'hE47;
		12'h5B4 : dout <= 12'hE45;
		12'h5B5 : dout <= 12'hE44;
		12'h5B6 : dout <= 12'hE42;
		12'h5B7 : dout <= 12'hE40;
		12'h5B8 : dout <= 12'hE3E;
		12'h5B9 : dout <= 12'hE3C;
		12'h5BA : dout <= 12'hE3A;
		12'h5BB : dout <= 12'hE38;
		12'h5BC : dout <= 12'hE36;
		12'h5BD : dout <= 12'hE34;
		12'h5BE : dout <= 12'hE32;
		12'h5BF : dout <= 12'hE30;
		12'h5C0 : dout <= 12'hE2E;
		12'h5C1 : dout <= 12'hE2C;
		12'h5C2 : dout <= 12'hE2A;
		12'h5C3 : dout <= 12'hE28;
		12'h5C4 : dout <= 12'hE26;
		12'h5C5 : dout <= 12'hE24;
		12'h5C6 : dout <= 12'hE22;
		12'h5C7 : dout <= 12'hE20;
		12'h5C8 : dout <= 12'hE1E;
		12'h5C9 : dout <= 12'hE1C;
		12'h5CA : dout <= 12'hE1A;
		12'h5CB : dout <= 12'hE18;
		12'h5CC : dout <= 12'hE16;
		12'h5CD : dout <= 12'hE14;
		12'h5CE : dout <= 12'hE12;
		12'h5CF : dout <= 12'hE10;
		12'h5D0 : dout <= 12'hE0E;
		12'h5D1 : dout <= 12'hE0B;
		12'h5D2 : dout <= 12'hE09;
		12'h5D3 : dout <= 12'hE07;
		12'h5D4 : dout <= 12'hE05;
		12'h5D5 : dout <= 12'hE03;
		12'h5D6 : dout <= 12'hE01;
		12'h5D7 : dout <= 12'hDFF;
		12'h5D8 : dout <= 12'hDFD;
		12'h5D9 : dout <= 12'hDFB;
		12'h5DA : dout <= 12'hDF9;
		12'h5DB : dout <= 12'hDF7;
		12'h5DC : dout <= 12'hDF5;
		12'h5DD : dout <= 12'hDF3;
		12'h5DE : dout <= 12'hDF0;
		12'h5DF : dout <= 12'hDEE;
		12'h5E0 : dout <= 12'hDEC;
		12'h5E1 : dout <= 12'hDEA;
		12'h5E2 : dout <= 12'hDE8;
		12'h5E3 : dout <= 12'hDE6;
		12'h5E4 : dout <= 12'hDE4;
		12'h5E5 : dout <= 12'hDE2;
		12'h5E6 : dout <= 12'hDE0;
		12'h5E7 : dout <= 12'hDDD;
		12'h5E8 : dout <= 12'hDDB;
		12'h5E9 : dout <= 12'hDD9;
		12'h5EA : dout <= 12'hDD7;
		12'h5EB : dout <= 12'hDD5;
		12'h5EC : dout <= 12'hDD3;
		12'h5ED : dout <= 12'hDD1;
		12'h5EE : dout <= 12'hDCE;
		12'h5EF : dout <= 12'hDCC;
		12'h5F0 : dout <= 12'hDCA;
		12'h5F1 : dout <= 12'hDC8;
		12'h5F2 : dout <= 12'hDC6;
		12'h5F3 : dout <= 12'hDC4;
		12'h5F4 : dout <= 12'hDC1;
		12'h5F5 : dout <= 12'hDBF;
		12'h5F6 : dout <= 12'hDBD;
		12'h5F7 : dout <= 12'hDBB;
		12'h5F8 : dout <= 12'hDB9;
		12'h5F9 : dout <= 12'hDB6;
		12'h5FA : dout <= 12'hDB4;
		12'h5FB : dout <= 12'hDB2;
		12'h5FC : dout <= 12'hDB0;
		12'h5FD : dout <= 12'hDAE;
		12'h5FE : dout <= 12'hDAB;
		12'h5FF : dout <= 12'hDA9;
		12'h600 : dout <= 12'hDA7;
		12'h601 : dout <= 12'hDA5;
		12'h602 : dout <= 12'hDA3;
		12'h603 : dout <= 12'hDA0;
		12'h604 : dout <= 12'hD9E;
		12'h605 : dout <= 12'hD9C;
		12'h606 : dout <= 12'hD9A;
		12'h607 : dout <= 12'hD97;
		12'h608 : dout <= 12'hD95;
		12'h609 : dout <= 12'hD93;
		12'h60A : dout <= 12'hD91;
		12'h60B : dout <= 12'hD8E;
		12'h60C : dout <= 12'hD8C;
		12'h60D : dout <= 12'hD8A;
		12'h60E : dout <= 12'hD88;
		12'h60F : dout <= 12'hD85;
		12'h610 : dout <= 12'hD83;
		12'h611 : dout <= 12'hD81;
		12'h612 : dout <= 12'hD7E;
		12'h613 : dout <= 12'hD7C;
		12'h614 : dout <= 12'hD7A;
		12'h615 : dout <= 12'hD78;
		12'h616 : dout <= 12'hD75;
		12'h617 : dout <= 12'hD73;
		12'h618 : dout <= 12'hD71;
		12'h619 : dout <= 12'hD6E;
		12'h61A : dout <= 12'hD6C;
		12'h61B : dout <= 12'hD6A;
		12'h61C : dout <= 12'hD67;
		12'h61D : dout <= 12'hD65;
		12'h61E : dout <= 12'hD63;
		12'h61F : dout <= 12'hD61;
		12'h620 : dout <= 12'hD5E;
		12'h621 : dout <= 12'hD5C;
		12'h622 : dout <= 12'hD5A;
		12'h623 : dout <= 12'hD57;
		12'h624 : dout <= 12'hD55;
		12'h625 : dout <= 12'hD53;
		12'h626 : dout <= 12'hD50;
		12'h627 : dout <= 12'hD4E;
		12'h628 : dout <= 12'hD4B;
		12'h629 : dout <= 12'hD49;
		12'h62A : dout <= 12'hD47;
		12'h62B : dout <= 12'hD44;
		12'h62C : dout <= 12'hD42;
		12'h62D : dout <= 12'hD40;
		12'h62E : dout <= 12'hD3D;
		12'h62F : dout <= 12'hD3B;
		12'h630 : dout <= 12'hD39;
		12'h631 : dout <= 12'hD36;
		12'h632 : dout <= 12'hD34;
		12'h633 : dout <= 12'hD31;
		12'h634 : dout <= 12'hD2F;
		12'h635 : dout <= 12'hD2D;
		12'h636 : dout <= 12'hD2A;
		12'h637 : dout <= 12'hD28;
		12'h638 : dout <= 12'hD25;
		12'h639 : dout <= 12'hD23;
		12'h63A : dout <= 12'hD21;
		12'h63B : dout <= 12'hD1E;
		12'h63C : dout <= 12'hD1C;
		12'h63D : dout <= 12'hD19;
		12'h63E : dout <= 12'hD17;
		12'h63F : dout <= 12'hD15;
		12'h640 : dout <= 12'hD12;
		12'h641 : dout <= 12'hD10;
		12'h642 : dout <= 12'hD0D;
		12'h643 : dout <= 12'hD0B;
		12'h644 : dout <= 12'hD08;
		12'h645 : dout <= 12'hD06;
		12'h646 : dout <= 12'hD03;
		12'h647 : dout <= 12'hD01;
		12'h648 : dout <= 12'hCFF;
		12'h649 : dout <= 12'hCFC;
		12'h64A : dout <= 12'hCFA;
		12'h64B : dout <= 12'hCF7;
		12'h64C : dout <= 12'hCF5;
		12'h64D : dout <= 12'hCF2;
		12'h64E : dout <= 12'hCF0;
		12'h64F : dout <= 12'hCED;
		12'h650 : dout <= 12'hCEB;
		12'h651 : dout <= 12'hCE8;
		12'h652 : dout <= 12'hCE6;
		12'h653 : dout <= 12'hCE3;
		12'h654 : dout <= 12'hCE1;
		12'h655 : dout <= 12'hCDE;
		12'h656 : dout <= 12'hCDC;
		12'h657 : dout <= 12'hCD9;
		12'h658 : dout <= 12'hCD7;
		12'h659 : dout <= 12'hCD4;
		12'h65A : dout <= 12'hCD2;
		12'h65B : dout <= 12'hCCF;
		12'h65C : dout <= 12'hCCD;
		12'h65D : dout <= 12'hCCA;
		12'h65E : dout <= 12'hCC8;
		12'h65F : dout <= 12'hCC5;
		12'h660 : dout <= 12'hCC3;
		12'h661 : dout <= 12'hCC0;
		12'h662 : dout <= 12'hCBE;
		12'h663 : dout <= 12'hCBB;
		12'h664 : dout <= 12'hCB9;
		12'h665 : dout <= 12'hCB6;
		12'h666 : dout <= 12'hCB4;
		12'h667 : dout <= 12'hCB1;
		12'h668 : dout <= 12'hCAF;
		12'h669 : dout <= 12'hCAC;
		12'h66A : dout <= 12'hCAA;
		12'h66B : dout <= 12'hCA7;
		12'h66C : dout <= 12'hCA4;
		12'h66D : dout <= 12'hCA2;
		12'h66E : dout <= 12'hC9F;
		12'h66F : dout <= 12'hC9D;
		12'h670 : dout <= 12'hC9A;
		12'h671 : dout <= 12'hC98;
		12'h672 : dout <= 12'hC95;
		12'h673 : dout <= 12'hC92;
		12'h674 : dout <= 12'hC90;
		12'h675 : dout <= 12'hC8D;
		12'h676 : dout <= 12'hC8B;
		12'h677 : dout <= 12'hC88;
		12'h678 : dout <= 12'hC86;
		12'h679 : dout <= 12'hC83;
		12'h67A : dout <= 12'hC80;
		12'h67B : dout <= 12'hC7E;
		12'h67C : dout <= 12'hC7B;
		12'h67D : dout <= 12'hC79;
		12'h67E : dout <= 12'hC76;
		12'h67F : dout <= 12'hC73;
		12'h680 : dout <= 12'hC71;
		12'h681 : dout <= 12'hC6E;
		12'h682 : dout <= 12'hC6C;
		12'h683 : dout <= 12'hC69;
		12'h684 : dout <= 12'hC66;
		12'h685 : dout <= 12'hC64;
		12'h686 : dout <= 12'hC61;
		12'h687 : dout <= 12'hC5E;
		12'h688 : dout <= 12'hC5C;
		12'h689 : dout <= 12'hC59;
		12'h68A : dout <= 12'hC57;
		12'h68B : dout <= 12'hC54;
		12'h68C : dout <= 12'hC51;
		12'h68D : dout <= 12'hC4F;
		12'h68E : dout <= 12'hC4C;
		12'h68F : dout <= 12'hC49;
		12'h690 : dout <= 12'hC47;
		12'h691 : dout <= 12'hC44;
		12'h692 : dout <= 12'hC41;
		12'h693 : dout <= 12'hC3F;
		12'h694 : dout <= 12'hC3C;
		12'h695 : dout <= 12'hC39;
		12'h696 : dout <= 12'hC37;
		12'h697 : dout <= 12'hC34;
		12'h698 : dout <= 12'hC31;
		12'h699 : dout <= 12'hC2F;
		12'h69A : dout <= 12'hC2C;
		12'h69B : dout <= 12'hC29;
		12'h69C : dout <= 12'hC27;
		12'h69D : dout <= 12'hC24;
		12'h69E : dout <= 12'hC21;
		12'h69F : dout <= 12'hC1F;
		12'h6A0 : dout <= 12'hC1C;
		12'h6A1 : dout <= 12'hC19;
		12'h6A2 : dout <= 12'hC16;
		12'h6A3 : dout <= 12'hC14;
		12'h6A4 : dout <= 12'hC11;
		12'h6A5 : dout <= 12'hC0E;
		12'h6A6 : dout <= 12'hC0C;
		12'h6A7 : dout <= 12'hC09;
		12'h6A8 : dout <= 12'hC06;
		12'h6A9 : dout <= 12'hC04;
		12'h6AA : dout <= 12'hC01;
		12'h6AB : dout <= 12'hBFE;
		12'h6AC : dout <= 12'hBFB;
		12'h6AD : dout <= 12'hBF9;
		12'h6AE : dout <= 12'hBF6;
		12'h6AF : dout <= 12'hBF3;
		12'h6B0 : dout <= 12'hBF0;
		12'h6B1 : dout <= 12'hBEE;
		12'h6B2 : dout <= 12'hBEB;
		12'h6B3 : dout <= 12'hBE8;
		12'h6B4 : dout <= 12'hBE6;
		12'h6B5 : dout <= 12'hBE3;
		12'h6B6 : dout <= 12'hBE0;
		12'h6B7 : dout <= 12'hBDD;
		12'h6B8 : dout <= 12'hBDB;
		12'h6B9 : dout <= 12'hBD8;
		12'h6BA : dout <= 12'hBD5;
		12'h6BB : dout <= 12'hBD2;
		12'h6BC : dout <= 12'hBD0;
		12'h6BD : dout <= 12'hBCD;
		12'h6BE : dout <= 12'hBCA;
		12'h6BF : dout <= 12'hBC7;
		12'h6C0 : dout <= 12'hBC4;
		12'h6C1 : dout <= 12'hBC2;
		12'h6C2 : dout <= 12'hBBF;
		12'h6C3 : dout <= 12'hBBC;
		12'h6C4 : dout <= 12'hBB9;
		12'h6C5 : dout <= 12'hBB7;
		12'h6C6 : dout <= 12'hBB4;
		12'h6C7 : dout <= 12'hBB1;
		12'h6C8 : dout <= 12'hBAE;
		12'h6C9 : dout <= 12'hBAB;
		12'h6CA : dout <= 12'hBA9;
		12'h6CB : dout <= 12'hBA6;
		12'h6CC : dout <= 12'hBA3;
		12'h6CD : dout <= 12'hBA0;
		12'h6CE : dout <= 12'hB9D;
		12'h6CF : dout <= 12'hB9B;
		12'h6D0 : dout <= 12'hB98;
		12'h6D1 : dout <= 12'hB95;
		12'h6D2 : dout <= 12'hB92;
		12'h6D3 : dout <= 12'hB8F;
		12'h6D4 : dout <= 12'hB8D;
		12'h6D5 : dout <= 12'hB8A;
		12'h6D6 : dout <= 12'hB87;
		12'h6D7 : dout <= 12'hB84;
		12'h6D8 : dout <= 12'hB81;
		12'h6D9 : dout <= 12'hB7F;
		12'h6DA : dout <= 12'hB7C;
		12'h6DB : dout <= 12'hB79;
		12'h6DC : dout <= 12'hB76;
		12'h6DD : dout <= 12'hB73;
		12'h6DE : dout <= 12'hB70;
		12'h6DF : dout <= 12'hB6E;
		12'h6E0 : dout <= 12'hB6B;
		12'h6E1 : dout <= 12'hB68;
		12'h6E2 : dout <= 12'hB65;
		12'h6E3 : dout <= 12'hB62;
		12'h6E4 : dout <= 12'hB5F;
		12'h6E5 : dout <= 12'hB5C;
		12'h6E6 : dout <= 12'hB5A;
		12'h6E7 : dout <= 12'hB57;
		12'h6E8 : dout <= 12'hB54;
		12'h6E9 : dout <= 12'hB51;
		12'h6EA : dout <= 12'hB4E;
		12'h6EB : dout <= 12'hB4B;
		12'h6EC : dout <= 12'hB48;
		12'h6ED : dout <= 12'hB46;
		12'h6EE : dout <= 12'hB43;
		12'h6EF : dout <= 12'hB40;
		12'h6F0 : dout <= 12'hB3D;
		12'h6F1 : dout <= 12'hB3A;
		12'h6F2 : dout <= 12'hB37;
		12'h6F3 : dout <= 12'hB34;
		12'h6F4 : dout <= 12'hB32;
		12'h6F5 : dout <= 12'hB2F;
		12'h6F6 : dout <= 12'hB2C;
		12'h6F7 : dout <= 12'hB29;
		12'h6F8 : dout <= 12'hB26;
		12'h6F9 : dout <= 12'hB23;
		12'h6FA : dout <= 12'hB20;
		12'h6FB : dout <= 12'hB1D;
		12'h6FC : dout <= 12'hB1A;
		12'h6FD : dout <= 12'hB18;
		12'h6FE : dout <= 12'hB15;
		12'h6FF : dout <= 12'hB12;
		12'h700 : dout <= 12'hB0F;
		12'h701 : dout <= 12'hB0C;
		12'h702 : dout <= 12'hB09;
		12'h703 : dout <= 12'hB06;
		12'h704 : dout <= 12'hB03;
		12'h705 : dout <= 12'hB00;
		12'h706 : dout <= 12'hAFD;
		12'h707 : dout <= 12'hAFB;
		12'h708 : dout <= 12'hAF8;
		12'h709 : dout <= 12'hAF5;
		12'h70A : dout <= 12'hAF2;
		12'h70B : dout <= 12'hAEF;
		12'h70C : dout <= 12'hAEC;
		12'h70D : dout <= 12'hAE9;
		12'h70E : dout <= 12'hAE6;
		12'h70F : dout <= 12'hAE3;
		12'h710 : dout <= 12'hAE0;
		12'h711 : dout <= 12'hADD;
		12'h712 : dout <= 12'hADA;
		12'h713 : dout <= 12'hAD7;
		12'h714 : dout <= 12'hAD4;
		12'h715 : dout <= 12'hAD2;
		12'h716 : dout <= 12'hACF;
		12'h717 : dout <= 12'hACC;
		12'h718 : dout <= 12'hAC9;
		12'h719 : dout <= 12'hAC6;
		12'h71A : dout <= 12'hAC3;
		12'h71B : dout <= 12'hAC0;
		12'h71C : dout <= 12'hABD;
		12'h71D : dout <= 12'hABA;
		12'h71E : dout <= 12'hAB7;
		12'h71F : dout <= 12'hAB4;
		12'h720 : dout <= 12'hAB1;
		12'h721 : dout <= 12'hAAE;
		12'h722 : dout <= 12'hAAB;
		12'h723 : dout <= 12'hAA8;
		12'h724 : dout <= 12'hAA5;
		12'h725 : dout <= 12'hAA2;
		12'h726 : dout <= 12'hA9F;
		12'h727 : dout <= 12'hA9C;
		12'h728 : dout <= 12'hA99;
		12'h729 : dout <= 12'hA96;
		12'h72A : dout <= 12'hA93;
		12'h72B : dout <= 12'hA90;
		12'h72C : dout <= 12'hA8E;
		12'h72D : dout <= 12'hA8B;
		12'h72E : dout <= 12'hA88;
		12'h72F : dout <= 12'hA85;
		12'h730 : dout <= 12'hA82;
		12'h731 : dout <= 12'hA7F;
		12'h732 : dout <= 12'hA7C;
		12'h733 : dout <= 12'hA79;
		12'h734 : dout <= 12'hA76;
		12'h735 : dout <= 12'hA73;
		12'h736 : dout <= 12'hA70;
		12'h737 : dout <= 12'hA6D;
		12'h738 : dout <= 12'hA6A;
		12'h739 : dout <= 12'hA67;
		12'h73A : dout <= 12'hA64;
		12'h73B : dout <= 12'hA61;
		12'h73C : dout <= 12'hA5E;
		12'h73D : dout <= 12'hA5B;
		12'h73E : dout <= 12'hA58;
		12'h73F : dout <= 12'hA55;
		12'h740 : dout <= 12'hA52;
		12'h741 : dout <= 12'hA4F;
		12'h742 : dout <= 12'hA4C;
		12'h743 : dout <= 12'hA49;
		12'h744 : dout <= 12'hA46;
		12'h745 : dout <= 12'hA43;
		12'h746 : dout <= 12'hA40;
		12'h747 : dout <= 12'hA3D;
		12'h748 : dout <= 12'hA3A;
		12'h749 : dout <= 12'hA37;
		12'h74A : dout <= 12'hA34;
		12'h74B : dout <= 12'hA31;
		12'h74C : dout <= 12'hA2E;
		12'h74D : dout <= 12'hA2B;
		12'h74E : dout <= 12'hA28;
		12'h74F : dout <= 12'hA24;
		12'h750 : dout <= 12'hA21;
		12'h751 : dout <= 12'hA1E;
		12'h752 : dout <= 12'hA1B;
		12'h753 : dout <= 12'hA18;
		12'h754 : dout <= 12'hA15;
		12'h755 : dout <= 12'hA12;
		12'h756 : dout <= 12'hA0F;
		12'h757 : dout <= 12'hA0C;
		12'h758 : dout <= 12'hA09;
		12'h759 : dout <= 12'hA06;
		12'h75A : dout <= 12'hA03;
		12'h75B : dout <= 12'hA00;
		12'h75C : dout <= 12'h9FD;
		12'h75D : dout <= 12'h9FA;
		12'h75E : dout <= 12'h9F7;
		12'h75F : dout <= 12'h9F4;
		12'h760 : dout <= 12'h9F1;
		12'h761 : dout <= 12'h9EE;
		12'h762 : dout <= 12'h9EB;
		12'h763 : dout <= 12'h9E8;
		12'h764 : dout <= 12'h9E5;
		12'h765 : dout <= 12'h9E2;
		12'h766 : dout <= 12'h9DF;
		12'h767 : dout <= 12'h9DC;
		12'h768 : dout <= 12'h9D8;
		12'h769 : dout <= 12'h9D5;
		12'h76A : dout <= 12'h9D2;
		12'h76B : dout <= 12'h9CF;
		12'h76C : dout <= 12'h9CC;
		12'h76D : dout <= 12'h9C9;
		12'h76E : dout <= 12'h9C6;
		12'h76F : dout <= 12'h9C3;
		12'h770 : dout <= 12'h9C0;
		12'h771 : dout <= 12'h9BD;
		12'h772 : dout <= 12'h9BA;
		12'h773 : dout <= 12'h9B7;
		12'h774 : dout <= 12'h9B4;
		12'h775 : dout <= 12'h9B1;
		12'h776 : dout <= 12'h9AE;
		12'h777 : dout <= 12'h9AB;
		12'h778 : dout <= 12'h9A7;
		12'h779 : dout <= 12'h9A4;
		12'h77A : dout <= 12'h9A1;
		12'h77B : dout <= 12'h99E;
		12'h77C : dout <= 12'h99B;
		12'h77D : dout <= 12'h998;
		12'h77E : dout <= 12'h995;
		12'h77F : dout <= 12'h992;
		12'h780 : dout <= 12'h98F;
		12'h781 : dout <= 12'h98C;
		12'h782 : dout <= 12'h989;
		12'h783 : dout <= 12'h986;
		12'h784 : dout <= 12'h983;
		12'h785 : dout <= 12'h97F;
		12'h786 : dout <= 12'h97C;
		12'h787 : dout <= 12'h979;
		12'h788 : dout <= 12'h976;
		12'h789 : dout <= 12'h973;
		12'h78A : dout <= 12'h970;
		12'h78B : dout <= 12'h96D;
		12'h78C : dout <= 12'h96A;
		12'h78D : dout <= 12'h967;
		12'h78E : dout <= 12'h964;
		12'h78F : dout <= 12'h961;
		12'h790 : dout <= 12'h95D;
		12'h791 : dout <= 12'h95A;
		12'h792 : dout <= 12'h957;
		12'h793 : dout <= 12'h954;
		12'h794 : dout <= 12'h951;
		12'h795 : dout <= 12'h94E;
		12'h796 : dout <= 12'h94B;
		12'h797 : dout <= 12'h948;
		12'h798 : dout <= 12'h945;
		12'h799 : dout <= 12'h942;
		12'h79A : dout <= 12'h93E;
		12'h79B : dout <= 12'h93B;
		12'h79C : dout <= 12'h938;
		12'h79D : dout <= 12'h935;
		12'h79E : dout <= 12'h932;
		12'h79F : dout <= 12'h92F;
		12'h7A0 : dout <= 12'h92C;
		12'h7A1 : dout <= 12'h929;
		12'h7A2 : dout <= 12'h926;
		12'h7A3 : dout <= 12'h923;
		12'h7A4 : dout <= 12'h91F;
		12'h7A5 : dout <= 12'h91C;
		12'h7A6 : dout <= 12'h919;
		12'h7A7 : dout <= 12'h916;
		12'h7A8 : dout <= 12'h913;
		12'h7A9 : dout <= 12'h910;
		12'h7AA : dout <= 12'h90D;
		12'h7AB : dout <= 12'h90A;
		12'h7AC : dout <= 12'h907;
		12'h7AD : dout <= 12'h903;
		12'h7AE : dout <= 12'h900;
		12'h7AF : dout <= 12'h8FD;
		12'h7B0 : dout <= 12'h8FA;
		12'h7B1 : dout <= 12'h8F7;
		12'h7B2 : dout <= 12'h8F4;
		12'h7B3 : dout <= 12'h8F1;
		12'h7B4 : dout <= 12'h8EE;
		12'h7B5 : dout <= 12'h8EA;
		12'h7B6 : dout <= 12'h8E7;
		12'h7B7 : dout <= 12'h8E4;
		12'h7B8 : dout <= 12'h8E1;
		12'h7B9 : dout <= 12'h8DE;
		12'h7BA : dout <= 12'h8DB;
		12'h7BB : dout <= 12'h8D8;
		12'h7BC : dout <= 12'h8D5;
		12'h7BD : dout <= 12'h8D2;
		12'h7BE : dout <= 12'h8CE;
		12'h7BF : dout <= 12'h8CB;
		12'h7C0 : dout <= 12'h8C8;
		12'h7C1 : dout <= 12'h8C5;
		12'h7C2 : dout <= 12'h8C2;
		12'h7C3 : dout <= 12'h8BF;
		12'h7C4 : dout <= 12'h8BC;
		12'h7C5 : dout <= 12'h8B9;
		12'h7C6 : dout <= 12'h8B5;
		12'h7C7 : dout <= 12'h8B2;
		12'h7C8 : dout <= 12'h8AF;
		12'h7C9 : dout <= 12'h8AC;
		12'h7CA : dout <= 12'h8A9;
		12'h7CB : dout <= 12'h8A6;
		12'h7CC : dout <= 12'h8A3;
		12'h7CD : dout <= 12'h89F;
		12'h7CE : dout <= 12'h89C;
		12'h7CF : dout <= 12'h899;
		12'h7D0 : dout <= 12'h896;
		12'h7D1 : dout <= 12'h893;
		12'h7D2 : dout <= 12'h890;
		12'h7D3 : dout <= 12'h88D;
		12'h7D4 : dout <= 12'h88A;
		12'h7D5 : dout <= 12'h886;
		12'h7D6 : dout <= 12'h883;
		12'h7D7 : dout <= 12'h880;
		12'h7D8 : dout <= 12'h87D;
		12'h7D9 : dout <= 12'h87A;
		12'h7DA : dout <= 12'h877;
		12'h7DB : dout <= 12'h874;
		12'h7DC : dout <= 12'h870;
		12'h7DD : dout <= 12'h86D;
		12'h7DE : dout <= 12'h86A;
		12'h7DF : dout <= 12'h867;
		12'h7E0 : dout <= 12'h864;
		12'h7E1 : dout <= 12'h861;
		12'h7E2 : dout <= 12'h85E;
		12'h7E3 : dout <= 12'h85B;
		12'h7E4 : dout <= 12'h857;
		12'h7E5 : dout <= 12'h854;
		12'h7E6 : dout <= 12'h851;
		12'h7E7 : dout <= 12'h84E;
		12'h7E8 : dout <= 12'h84B;
		12'h7E9 : dout <= 12'h848;
		12'h7EA : dout <= 12'h845;
		12'h7EB : dout <= 12'h841;
		12'h7EC : dout <= 12'h83E;
		12'h7ED : dout <= 12'h83B;
		12'h7EE : dout <= 12'h838;
		12'h7EF : dout <= 12'h835;
		12'h7F0 : dout <= 12'h832;
		12'h7F1 : dout <= 12'h82F;
		12'h7F2 : dout <= 12'h82B;
		12'h7F3 : dout <= 12'h828;
		12'h7F4 : dout <= 12'h825;
		12'h7F5 : dout <= 12'h822;
		12'h7F6 : dout <= 12'h81F;
		12'h7F7 : dout <= 12'h81C;
		12'h7F8 : dout <= 12'h819;
		12'h7F9 : dout <= 12'h815;
		12'h7FA : dout <= 12'h812;
		12'h7FB : dout <= 12'h80F;
		12'h7FC : dout <= 12'h80C;
		12'h7FD : dout <= 12'h809;
		12'h7FE : dout <= 12'h806;
		12'h7FF : dout <= 12'h803;
		12'h800 : dout <= 12'h800;
		12'h801 : dout <= 12'h7FC;
		12'h802 : dout <= 12'h7F9;
		12'h803 : dout <= 12'h7F6;
		12'h804 : dout <= 12'h7F3;
		12'h805 : dout <= 12'h7F0;
		12'h806 : dout <= 12'h7ED;
		12'h807 : dout <= 12'h7EA;
		12'h808 : dout <= 12'h7E6;
		12'h809 : dout <= 12'h7E3;
		12'h80A : dout <= 12'h7E0;
		12'h80B : dout <= 12'h7DD;
		12'h80C : dout <= 12'h7DA;
		12'h80D : dout <= 12'h7D7;
		12'h80E : dout <= 12'h7D4;
		12'h80F : dout <= 12'h7D0;
		12'h810 : dout <= 12'h7CD;
		12'h811 : dout <= 12'h7CA;
		12'h812 : dout <= 12'h7C7;
		12'h813 : dout <= 12'h7C4;
		12'h814 : dout <= 12'h7C1;
		12'h815 : dout <= 12'h7BE;
		12'h816 : dout <= 12'h7BA;
		12'h817 : dout <= 12'h7B7;
		12'h818 : dout <= 12'h7B4;
		12'h819 : dout <= 12'h7B1;
		12'h81A : dout <= 12'h7AE;
		12'h81B : dout <= 12'h7AB;
		12'h81C : dout <= 12'h7A8;
		12'h81D : dout <= 12'h7A4;
		12'h81E : dout <= 12'h7A1;
		12'h81F : dout <= 12'h79E;
		12'h820 : dout <= 12'h79B;
		12'h821 : dout <= 12'h798;
		12'h822 : dout <= 12'h795;
		12'h823 : dout <= 12'h792;
		12'h824 : dout <= 12'h78F;
		12'h825 : dout <= 12'h78B;
		12'h826 : dout <= 12'h788;
		12'h827 : dout <= 12'h785;
		12'h828 : dout <= 12'h782;
		12'h829 : dout <= 12'h77F;
		12'h82A : dout <= 12'h77C;
		12'h82B : dout <= 12'h779;
		12'h82C : dout <= 12'h775;
		12'h82D : dout <= 12'h772;
		12'h82E : dout <= 12'h76F;
		12'h82F : dout <= 12'h76C;
		12'h830 : dout <= 12'h769;
		12'h831 : dout <= 12'h766;
		12'h832 : dout <= 12'h763;
		12'h833 : dout <= 12'h760;
		12'h834 : dout <= 12'h75C;
		12'h835 : dout <= 12'h759;
		12'h836 : dout <= 12'h756;
		12'h837 : dout <= 12'h753;
		12'h838 : dout <= 12'h750;
		12'h839 : dout <= 12'h74D;
		12'h83A : dout <= 12'h74A;
		12'h83B : dout <= 12'h746;
		12'h83C : dout <= 12'h743;
		12'h83D : dout <= 12'h740;
		12'h83E : dout <= 12'h73D;
		12'h83F : dout <= 12'h73A;
		12'h840 : dout <= 12'h737;
		12'h841 : dout <= 12'h734;
		12'h842 : dout <= 12'h731;
		12'h843 : dout <= 12'h72D;
		12'h844 : dout <= 12'h72A;
		12'h845 : dout <= 12'h727;
		12'h846 : dout <= 12'h724;
		12'h847 : dout <= 12'h721;
		12'h848 : dout <= 12'h71E;
		12'h849 : dout <= 12'h71B;
		12'h84A : dout <= 12'h718;
		12'h84B : dout <= 12'h715;
		12'h84C : dout <= 12'h711;
		12'h84D : dout <= 12'h70E;
		12'h84E : dout <= 12'h70B;
		12'h84F : dout <= 12'h708;
		12'h850 : dout <= 12'h705;
		12'h851 : dout <= 12'h702;
		12'h852 : dout <= 12'h6FF;
		12'h853 : dout <= 12'h6FC;
		12'h854 : dout <= 12'h6F8;
		12'h855 : dout <= 12'h6F5;
		12'h856 : dout <= 12'h6F2;
		12'h857 : dout <= 12'h6EF;
		12'h858 : dout <= 12'h6EC;
		12'h859 : dout <= 12'h6E9;
		12'h85A : dout <= 12'h6E6;
		12'h85B : dout <= 12'h6E3;
		12'h85C : dout <= 12'h6E0;
		12'h85D : dout <= 12'h6DC;
		12'h85E : dout <= 12'h6D9;
		12'h85F : dout <= 12'h6D6;
		12'h860 : dout <= 12'h6D3;
		12'h861 : dout <= 12'h6D0;
		12'h862 : dout <= 12'h6CD;
		12'h863 : dout <= 12'h6CA;
		12'h864 : dout <= 12'h6C7;
		12'h865 : dout <= 12'h6C4;
		12'h866 : dout <= 12'h6C1;
		12'h867 : dout <= 12'h6BD;
		12'h868 : dout <= 12'h6BA;
		12'h869 : dout <= 12'h6B7;
		12'h86A : dout <= 12'h6B4;
		12'h86B : dout <= 12'h6B1;
		12'h86C : dout <= 12'h6AE;
		12'h86D : dout <= 12'h6AB;
		12'h86E : dout <= 12'h6A8;
		12'h86F : dout <= 12'h6A5;
		12'h870 : dout <= 12'h6A2;
		12'h871 : dout <= 12'h69E;
		12'h872 : dout <= 12'h69B;
		12'h873 : dout <= 12'h698;
		12'h874 : dout <= 12'h695;
		12'h875 : dout <= 12'h692;
		12'h876 : dout <= 12'h68F;
		12'h877 : dout <= 12'h68C;
		12'h878 : dout <= 12'h689;
		12'h879 : dout <= 12'h686;
		12'h87A : dout <= 12'h683;
		12'h87B : dout <= 12'h680;
		12'h87C : dout <= 12'h67C;
		12'h87D : dout <= 12'h679;
		12'h87E : dout <= 12'h676;
		12'h87F : dout <= 12'h673;
		12'h880 : dout <= 12'h670;
		12'h881 : dout <= 12'h66D;
		12'h882 : dout <= 12'h66A;
		12'h883 : dout <= 12'h667;
		12'h884 : dout <= 12'h664;
		12'h885 : dout <= 12'h661;
		12'h886 : dout <= 12'h65E;
		12'h887 : dout <= 12'h65B;
		12'h888 : dout <= 12'h658;
		12'h889 : dout <= 12'h654;
		12'h88A : dout <= 12'h651;
		12'h88B : dout <= 12'h64E;
		12'h88C : dout <= 12'h64B;
		12'h88D : dout <= 12'h648;
		12'h88E : dout <= 12'h645;
		12'h88F : dout <= 12'h642;
		12'h890 : dout <= 12'h63F;
		12'h891 : dout <= 12'h63C;
		12'h892 : dout <= 12'h639;
		12'h893 : dout <= 12'h636;
		12'h894 : dout <= 12'h633;
		12'h895 : dout <= 12'h630;
		12'h896 : dout <= 12'h62D;
		12'h897 : dout <= 12'h62A;
		12'h898 : dout <= 12'h627;
		12'h899 : dout <= 12'h623;
		12'h89A : dout <= 12'h620;
		12'h89B : dout <= 12'h61D;
		12'h89C : dout <= 12'h61A;
		12'h89D : dout <= 12'h617;
		12'h89E : dout <= 12'h614;
		12'h89F : dout <= 12'h611;
		12'h8A0 : dout <= 12'h60E;
		12'h8A1 : dout <= 12'h60B;
		12'h8A2 : dout <= 12'h608;
		12'h8A3 : dout <= 12'h605;
		12'h8A4 : dout <= 12'h602;
		12'h8A5 : dout <= 12'h5FF;
		12'h8A6 : dout <= 12'h5FC;
		12'h8A7 : dout <= 12'h5F9;
		12'h8A8 : dout <= 12'h5F6;
		12'h8A9 : dout <= 12'h5F3;
		12'h8AA : dout <= 12'h5F0;
		12'h8AB : dout <= 12'h5ED;
		12'h8AC : dout <= 12'h5EA;
		12'h8AD : dout <= 12'h5E7;
		12'h8AE : dout <= 12'h5E4;
		12'h8AF : dout <= 12'h5E1;
		12'h8B0 : dout <= 12'h5DE;
		12'h8B1 : dout <= 12'h5DB;
		12'h8B2 : dout <= 12'h5D7;
		12'h8B3 : dout <= 12'h5D4;
		12'h8B4 : dout <= 12'h5D1;
		12'h8B5 : dout <= 12'h5CE;
		12'h8B6 : dout <= 12'h5CB;
		12'h8B7 : dout <= 12'h5C8;
		12'h8B8 : dout <= 12'h5C5;
		12'h8B9 : dout <= 12'h5C2;
		12'h8BA : dout <= 12'h5BF;
		12'h8BB : dout <= 12'h5BC;
		12'h8BC : dout <= 12'h5B9;
		12'h8BD : dout <= 12'h5B6;
		12'h8BE : dout <= 12'h5B3;
		12'h8BF : dout <= 12'h5B0;
		12'h8C0 : dout <= 12'h5AD;
		12'h8C1 : dout <= 12'h5AA;
		12'h8C2 : dout <= 12'h5A7;
		12'h8C3 : dout <= 12'h5A4;
		12'h8C4 : dout <= 12'h5A1;
		12'h8C5 : dout <= 12'h59E;
		12'h8C6 : dout <= 12'h59B;
		12'h8C7 : dout <= 12'h598;
		12'h8C8 : dout <= 12'h595;
		12'h8C9 : dout <= 12'h592;
		12'h8CA : dout <= 12'h58F;
		12'h8CB : dout <= 12'h58C;
		12'h8CC : dout <= 12'h589;
		12'h8CD : dout <= 12'h586;
		12'h8CE : dout <= 12'h583;
		12'h8CF : dout <= 12'h580;
		12'h8D0 : dout <= 12'h57D;
		12'h8D1 : dout <= 12'h57A;
		12'h8D2 : dout <= 12'h577;
		12'h8D3 : dout <= 12'h574;
		12'h8D4 : dout <= 12'h571;
		12'h8D5 : dout <= 12'h56F;
		12'h8D6 : dout <= 12'h56C;
		12'h8D7 : dout <= 12'h569;
		12'h8D8 : dout <= 12'h566;
		12'h8D9 : dout <= 12'h563;
		12'h8DA : dout <= 12'h560;
		12'h8DB : dout <= 12'h55D;
		12'h8DC : dout <= 12'h55A;
		12'h8DD : dout <= 12'h557;
		12'h8DE : dout <= 12'h554;
		12'h8DF : dout <= 12'h551;
		12'h8E0 : dout <= 12'h54E;
		12'h8E1 : dout <= 12'h54B;
		12'h8E2 : dout <= 12'h548;
		12'h8E3 : dout <= 12'h545;
		12'h8E4 : dout <= 12'h542;
		12'h8E5 : dout <= 12'h53F;
		12'h8E6 : dout <= 12'h53C;
		12'h8E7 : dout <= 12'h539;
		12'h8E8 : dout <= 12'h536;
		12'h8E9 : dout <= 12'h533;
		12'h8EA : dout <= 12'h530;
		12'h8EB : dout <= 12'h52D;
		12'h8EC : dout <= 12'h52B;
		12'h8ED : dout <= 12'h528;
		12'h8EE : dout <= 12'h525;
		12'h8EF : dout <= 12'h522;
		12'h8F0 : dout <= 12'h51F;
		12'h8F1 : dout <= 12'h51C;
		12'h8F2 : dout <= 12'h519;
		12'h8F3 : dout <= 12'h516;
		12'h8F4 : dout <= 12'h513;
		12'h8F5 : dout <= 12'h510;
		12'h8F6 : dout <= 12'h50D;
		12'h8F7 : dout <= 12'h50A;
		12'h8F8 : dout <= 12'h507;
		12'h8F9 : dout <= 12'h504;
		12'h8FA : dout <= 12'h502;
		12'h8FB : dout <= 12'h4FF;
		12'h8FC : dout <= 12'h4FC;
		12'h8FD : dout <= 12'h4F9;
		12'h8FE : dout <= 12'h4F6;
		12'h8FF : dout <= 12'h4F3;
		12'h900 : dout <= 12'h4F0;
		12'h901 : dout <= 12'h4ED;
		12'h902 : dout <= 12'h4EA;
		12'h903 : dout <= 12'h4E7;
		12'h904 : dout <= 12'h4E5;
		12'h905 : dout <= 12'h4E2;
		12'h906 : dout <= 12'h4DF;
		12'h907 : dout <= 12'h4DC;
		12'h908 : dout <= 12'h4D9;
		12'h909 : dout <= 12'h4D6;
		12'h90A : dout <= 12'h4D3;
		12'h90B : dout <= 12'h4D0;
		12'h90C : dout <= 12'h4CD;
		12'h90D : dout <= 12'h4CB;
		12'h90E : dout <= 12'h4C8;
		12'h90F : dout <= 12'h4C5;
		12'h910 : dout <= 12'h4C2;
		12'h911 : dout <= 12'h4BF;
		12'h912 : dout <= 12'h4BC;
		12'h913 : dout <= 12'h4B9;
		12'h914 : dout <= 12'h4B7;
		12'h915 : dout <= 12'h4B4;
		12'h916 : dout <= 12'h4B1;
		12'h917 : dout <= 12'h4AE;
		12'h918 : dout <= 12'h4AB;
		12'h919 : dout <= 12'h4A8;
		12'h91A : dout <= 12'h4A5;
		12'h91B : dout <= 12'h4A3;
		12'h91C : dout <= 12'h4A0;
		12'h91D : dout <= 12'h49D;
		12'h91E : dout <= 12'h49A;
		12'h91F : dout <= 12'h497;
		12'h920 : dout <= 12'h494;
		12'h921 : dout <= 12'h491;
		12'h922 : dout <= 12'h48F;
		12'h923 : dout <= 12'h48C;
		12'h924 : dout <= 12'h489;
		12'h925 : dout <= 12'h486;
		12'h926 : dout <= 12'h483;
		12'h927 : dout <= 12'h480;
		12'h928 : dout <= 12'h47E;
		12'h929 : dout <= 12'h47B;
		12'h92A : dout <= 12'h478;
		12'h92B : dout <= 12'h475;
		12'h92C : dout <= 12'h472;
		12'h92D : dout <= 12'h470;
		12'h92E : dout <= 12'h46D;
		12'h92F : dout <= 12'h46A;
		12'h930 : dout <= 12'h467;
		12'h931 : dout <= 12'h464;
		12'h932 : dout <= 12'h462;
		12'h933 : dout <= 12'h45F;
		12'h934 : dout <= 12'h45C;
		12'h935 : dout <= 12'h459;
		12'h936 : dout <= 12'h456;
		12'h937 : dout <= 12'h454;
		12'h938 : dout <= 12'h451;
		12'h939 : dout <= 12'h44E;
		12'h93A : dout <= 12'h44B;
		12'h93B : dout <= 12'h448;
		12'h93C : dout <= 12'h446;
		12'h93D : dout <= 12'h443;
		12'h93E : dout <= 12'h440;
		12'h93F : dout <= 12'h43D;
		12'h940 : dout <= 12'h43B;
		12'h941 : dout <= 12'h438;
		12'h942 : dout <= 12'h435;
		12'h943 : dout <= 12'h432;
		12'h944 : dout <= 12'h42F;
		12'h945 : dout <= 12'h42D;
		12'h946 : dout <= 12'h42A;
		12'h947 : dout <= 12'h427;
		12'h948 : dout <= 12'h424;
		12'h949 : dout <= 12'h422;
		12'h94A : dout <= 12'h41F;
		12'h94B : dout <= 12'h41C;
		12'h94C : dout <= 12'h419;
		12'h94D : dout <= 12'h417;
		12'h94E : dout <= 12'h414;
		12'h94F : dout <= 12'h411;
		12'h950 : dout <= 12'h40F;
		12'h951 : dout <= 12'h40C;
		12'h952 : dout <= 12'h409;
		12'h953 : dout <= 12'h406;
		12'h954 : dout <= 12'h404;
		12'h955 : dout <= 12'h401;
		12'h956 : dout <= 12'h3FE;
		12'h957 : dout <= 12'h3FB;
		12'h958 : dout <= 12'h3F9;
		12'h959 : dout <= 12'h3F6;
		12'h95A : dout <= 12'h3F3;
		12'h95B : dout <= 12'h3F1;
		12'h95C : dout <= 12'h3EE;
		12'h95D : dout <= 12'h3EB;
		12'h95E : dout <= 12'h3E9;
		12'h95F : dout <= 12'h3E6;
		12'h960 : dout <= 12'h3E3;
		12'h961 : dout <= 12'h3E0;
		12'h962 : dout <= 12'h3DE;
		12'h963 : dout <= 12'h3DB;
		12'h964 : dout <= 12'h3D8;
		12'h965 : dout <= 12'h3D6;
		12'h966 : dout <= 12'h3D3;
		12'h967 : dout <= 12'h3D0;
		12'h968 : dout <= 12'h3CE;
		12'h969 : dout <= 12'h3CB;
		12'h96A : dout <= 12'h3C8;
		12'h96B : dout <= 12'h3C6;
		12'h96C : dout <= 12'h3C3;
		12'h96D : dout <= 12'h3C0;
		12'h96E : dout <= 12'h3BE;
		12'h96F : dout <= 12'h3BB;
		12'h970 : dout <= 12'h3B8;
		12'h971 : dout <= 12'h3B6;
		12'h972 : dout <= 12'h3B3;
		12'h973 : dout <= 12'h3B0;
		12'h974 : dout <= 12'h3AE;
		12'h975 : dout <= 12'h3AB;
		12'h976 : dout <= 12'h3A8;
		12'h977 : dout <= 12'h3A6;
		12'h978 : dout <= 12'h3A3;
		12'h979 : dout <= 12'h3A1;
		12'h97A : dout <= 12'h39E;
		12'h97B : dout <= 12'h39B;
		12'h97C : dout <= 12'h399;
		12'h97D : dout <= 12'h396;
		12'h97E : dout <= 12'h393;
		12'h97F : dout <= 12'h391;
		12'h980 : dout <= 12'h38E;
		12'h981 : dout <= 12'h38C;
		12'h982 : dout <= 12'h389;
		12'h983 : dout <= 12'h386;
		12'h984 : dout <= 12'h384;
		12'h985 : dout <= 12'h381;
		12'h986 : dout <= 12'h37F;
		12'h987 : dout <= 12'h37C;
		12'h988 : dout <= 12'h379;
		12'h989 : dout <= 12'h377;
		12'h98A : dout <= 12'h374;
		12'h98B : dout <= 12'h372;
		12'h98C : dout <= 12'h36F;
		12'h98D : dout <= 12'h36D;
		12'h98E : dout <= 12'h36A;
		12'h98F : dout <= 12'h367;
		12'h990 : dout <= 12'h365;
		12'h991 : dout <= 12'h362;
		12'h992 : dout <= 12'h360;
		12'h993 : dout <= 12'h35D;
		12'h994 : dout <= 12'h35B;
		12'h995 : dout <= 12'h358;
		12'h996 : dout <= 12'h355;
		12'h997 : dout <= 12'h353;
		12'h998 : dout <= 12'h350;
		12'h999 : dout <= 12'h34E;
		12'h99A : dout <= 12'h34B;
		12'h99B : dout <= 12'h349;
		12'h99C : dout <= 12'h346;
		12'h99D : dout <= 12'h344;
		12'h99E : dout <= 12'h341;
		12'h99F : dout <= 12'h33F;
		12'h9A0 : dout <= 12'h33C;
		12'h9A1 : dout <= 12'h33A;
		12'h9A2 : dout <= 12'h337;
		12'h9A3 : dout <= 12'h335;
		12'h9A4 : dout <= 12'h332;
		12'h9A5 : dout <= 12'h330;
		12'h9A6 : dout <= 12'h32D;
		12'h9A7 : dout <= 12'h32B;
		12'h9A8 : dout <= 12'h328;
		12'h9A9 : dout <= 12'h326;
		12'h9AA : dout <= 12'h323;
		12'h9AB : dout <= 12'h321;
		12'h9AC : dout <= 12'h31E;
		12'h9AD : dout <= 12'h31C;
		12'h9AE : dout <= 12'h319;
		12'h9AF : dout <= 12'h317;
		12'h9B0 : dout <= 12'h314;
		12'h9B1 : dout <= 12'h312;
		12'h9B2 : dout <= 12'h30F;
		12'h9B3 : dout <= 12'h30D;
		12'h9B4 : dout <= 12'h30A;
		12'h9B5 : dout <= 12'h308;
		12'h9B6 : dout <= 12'h305;
		12'h9B7 : dout <= 12'h303;
		12'h9B8 : dout <= 12'h300;
		12'h9B9 : dout <= 12'h2FE;
		12'h9BA : dout <= 12'h2FC;
		12'h9BB : dout <= 12'h2F9;
		12'h9BC : dout <= 12'h2F7;
		12'h9BD : dout <= 12'h2F4;
		12'h9BE : dout <= 12'h2F2;
		12'h9BF : dout <= 12'h2EF;
		12'h9C0 : dout <= 12'h2ED;
		12'h9C1 : dout <= 12'h2EA;
		12'h9C2 : dout <= 12'h2E8;
		12'h9C3 : dout <= 12'h2E6;
		12'h9C4 : dout <= 12'h2E3;
		12'h9C5 : dout <= 12'h2E1;
		12'h9C6 : dout <= 12'h2DE;
		12'h9C7 : dout <= 12'h2DC;
		12'h9C8 : dout <= 12'h2DA;
		12'h9C9 : dout <= 12'h2D7;
		12'h9CA : dout <= 12'h2D5;
		12'h9CB : dout <= 12'h2D2;
		12'h9CC : dout <= 12'h2D0;
		12'h9CD : dout <= 12'h2CE;
		12'h9CE : dout <= 12'h2CB;
		12'h9CF : dout <= 12'h2C9;
		12'h9D0 : dout <= 12'h2C6;
		12'h9D1 : dout <= 12'h2C4;
		12'h9D2 : dout <= 12'h2C2;
		12'h9D3 : dout <= 12'h2BF;
		12'h9D4 : dout <= 12'h2BD;
		12'h9D5 : dout <= 12'h2BB;
		12'h9D6 : dout <= 12'h2B8;
		12'h9D7 : dout <= 12'h2B6;
		12'h9D8 : dout <= 12'h2B4;
		12'h9D9 : dout <= 12'h2B1;
		12'h9DA : dout <= 12'h2AF;
		12'h9DB : dout <= 12'h2AC;
		12'h9DC : dout <= 12'h2AA;
		12'h9DD : dout <= 12'h2A8;
		12'h9DE : dout <= 12'h2A5;
		12'h9DF : dout <= 12'h2A3;
		12'h9E0 : dout <= 12'h2A1;
		12'h9E1 : dout <= 12'h29E;
		12'h9E2 : dout <= 12'h29C;
		12'h9E3 : dout <= 12'h29A;
		12'h9E4 : dout <= 12'h298;
		12'h9E5 : dout <= 12'h295;
		12'h9E6 : dout <= 12'h293;
		12'h9E7 : dout <= 12'h291;
		12'h9E8 : dout <= 12'h28E;
		12'h9E9 : dout <= 12'h28C;
		12'h9EA : dout <= 12'h28A;
		12'h9EB : dout <= 12'h287;
		12'h9EC : dout <= 12'h285;
		12'h9ED : dout <= 12'h283;
		12'h9EE : dout <= 12'h281;
		12'h9EF : dout <= 12'h27E;
		12'h9F0 : dout <= 12'h27C;
		12'h9F1 : dout <= 12'h27A;
		12'h9F2 : dout <= 12'h277;
		12'h9F3 : dout <= 12'h275;
		12'h9F4 : dout <= 12'h273;
		12'h9F5 : dout <= 12'h271;
		12'h9F6 : dout <= 12'h26E;
		12'h9F7 : dout <= 12'h26C;
		12'h9F8 : dout <= 12'h26A;
		12'h9F9 : dout <= 12'h268;
		12'h9FA : dout <= 12'h265;
		12'h9FB : dout <= 12'h263;
		12'h9FC : dout <= 12'h261;
		12'h9FD : dout <= 12'h25F;
		12'h9FE : dout <= 12'h25C;
		12'h9FF : dout <= 12'h25A;
		12'hA00 : dout <= 12'h258;
		12'hA01 : dout <= 12'h256;
		12'hA02 : dout <= 12'h254;
		12'hA03 : dout <= 12'h251;
		12'hA04 : dout <= 12'h24F;
		12'hA05 : dout <= 12'h24D;
		12'hA06 : dout <= 12'h24B;
		12'hA07 : dout <= 12'h249;
		12'hA08 : dout <= 12'h246;
		12'hA09 : dout <= 12'h244;
		12'hA0A : dout <= 12'h242;
		12'hA0B : dout <= 12'h240;
		12'hA0C : dout <= 12'h23E;
		12'hA0D : dout <= 12'h23B;
		12'hA0E : dout <= 12'h239;
		12'hA0F : dout <= 12'h237;
		12'hA10 : dout <= 12'h235;
		12'hA11 : dout <= 12'h233;
		12'hA12 : dout <= 12'h231;
		12'hA13 : dout <= 12'h22E;
		12'hA14 : dout <= 12'h22C;
		12'hA15 : dout <= 12'h22A;
		12'hA16 : dout <= 12'h228;
		12'hA17 : dout <= 12'h226;
		12'hA18 : dout <= 12'h224;
		12'hA19 : dout <= 12'h222;
		12'hA1A : dout <= 12'h21F;
		12'hA1B : dout <= 12'h21D;
		12'hA1C : dout <= 12'h21B;
		12'hA1D : dout <= 12'h219;
		12'hA1E : dout <= 12'h217;
		12'hA1F : dout <= 12'h215;
		12'hA20 : dout <= 12'h213;
		12'hA21 : dout <= 12'h211;
		12'hA22 : dout <= 12'h20F;
		12'hA23 : dout <= 12'h20C;
		12'hA24 : dout <= 12'h20A;
		12'hA25 : dout <= 12'h208;
		12'hA26 : dout <= 12'h206;
		12'hA27 : dout <= 12'h204;
		12'hA28 : dout <= 12'h202;
		12'hA29 : dout <= 12'h200;
		12'hA2A : dout <= 12'h1FE;
		12'hA2B : dout <= 12'h1FC;
		12'hA2C : dout <= 12'h1FA;
		12'hA2D : dout <= 12'h1F8;
		12'hA2E : dout <= 12'h1F6;
		12'hA2F : dout <= 12'h1F4;
		12'hA30 : dout <= 12'h1F1;
		12'hA31 : dout <= 12'h1EF;
		12'hA32 : dout <= 12'h1ED;
		12'hA33 : dout <= 12'h1EB;
		12'hA34 : dout <= 12'h1E9;
		12'hA35 : dout <= 12'h1E7;
		12'hA36 : dout <= 12'h1E5;
		12'hA37 : dout <= 12'h1E3;
		12'hA38 : dout <= 12'h1E1;
		12'hA39 : dout <= 12'h1DF;
		12'hA3A : dout <= 12'h1DD;
		12'hA3B : dout <= 12'h1DB;
		12'hA3C : dout <= 12'h1D9;
		12'hA3D : dout <= 12'h1D7;
		12'hA3E : dout <= 12'h1D5;
		12'hA3F : dout <= 12'h1D3;
		12'hA40 : dout <= 12'h1D1;
		12'hA41 : dout <= 12'h1CF;
		12'hA42 : dout <= 12'h1CD;
		12'hA43 : dout <= 12'h1CB;
		12'hA44 : dout <= 12'h1C9;
		12'hA45 : dout <= 12'h1C7;
		12'hA46 : dout <= 12'h1C5;
		12'hA47 : dout <= 12'h1C3;
		12'hA48 : dout <= 12'h1C1;
		12'hA49 : dout <= 12'h1BF;
		12'hA4A : dout <= 12'h1BD;
		12'hA4B : dout <= 12'h1BB;
		12'hA4C : dout <= 12'h1BA;
		12'hA4D : dout <= 12'h1B8;
		12'hA4E : dout <= 12'h1B6;
		12'hA4F : dout <= 12'h1B4;
		12'hA50 : dout <= 12'h1B2;
		12'hA51 : dout <= 12'h1B0;
		12'hA52 : dout <= 12'h1AE;
		12'hA53 : dout <= 12'h1AC;
		12'hA54 : dout <= 12'h1AA;
		12'hA55 : dout <= 12'h1A8;
		12'hA56 : dout <= 12'h1A6;
		12'hA57 : dout <= 12'h1A4;
		12'hA58 : dout <= 12'h1A2;
		12'hA59 : dout <= 12'h1A1;
		12'hA5A : dout <= 12'h19F;
		12'hA5B : dout <= 12'h19D;
		12'hA5C : dout <= 12'h19B;
		12'hA5D : dout <= 12'h199;
		12'hA5E : dout <= 12'h197;
		12'hA5F : dout <= 12'h195;
		12'hA60 : dout <= 12'h193;
		12'hA61 : dout <= 12'h191;
		12'hA62 : dout <= 12'h190;
		12'hA63 : dout <= 12'h18E;
		12'hA64 : dout <= 12'h18C;
		12'hA65 : dout <= 12'h18A;
		12'hA66 : dout <= 12'h188;
		12'hA67 : dout <= 12'h186;
		12'hA68 : dout <= 12'h184;
		12'hA69 : dout <= 12'h183;
		12'hA6A : dout <= 12'h181;
		12'hA6B : dout <= 12'h17F;
		12'hA6C : dout <= 12'h17D;
		12'hA6D : dout <= 12'h17B;
		12'hA6E : dout <= 12'h17A;
		12'hA6F : dout <= 12'h178;
		12'hA70 : dout <= 12'h176;
		12'hA71 : dout <= 12'h174;
		12'hA72 : dout <= 12'h172;
		12'hA73 : dout <= 12'h170;
		12'hA74 : dout <= 12'h16F;
		12'hA75 : dout <= 12'h16D;
		12'hA76 : dout <= 12'h16B;
		12'hA77 : dout <= 12'h169;
		12'hA78 : dout <= 12'h168;
		12'hA79 : dout <= 12'h166;
		12'hA7A : dout <= 12'h164;
		12'hA7B : dout <= 12'h162;
		12'hA7C : dout <= 12'h160;
		12'hA7D : dout <= 12'h15F;
		12'hA7E : dout <= 12'h15D;
		12'hA7F : dout <= 12'h15B;
		12'hA80 : dout <= 12'h159;
		12'hA81 : dout <= 12'h158;
		12'hA82 : dout <= 12'h156;
		12'hA83 : dout <= 12'h154;
		12'hA84 : dout <= 12'h153;
		12'hA85 : dout <= 12'h151;
		12'hA86 : dout <= 12'h14F;
		12'hA87 : dout <= 12'h14D;
		12'hA88 : dout <= 12'h14C;
		12'hA89 : dout <= 12'h14A;
		12'hA8A : dout <= 12'h148;
		12'hA8B : dout <= 12'h147;
		12'hA8C : dout <= 12'h145;
		12'hA8D : dout <= 12'h143;
		12'hA8E : dout <= 12'h141;
		12'hA8F : dout <= 12'h140;
		12'hA90 : dout <= 12'h13E;
		12'hA91 : dout <= 12'h13C;
		12'hA92 : dout <= 12'h13B;
		12'hA93 : dout <= 12'h139;
		12'hA94 : dout <= 12'h137;
		12'hA95 : dout <= 12'h136;
		12'hA96 : dout <= 12'h134;
		12'hA97 : dout <= 12'h132;
		12'hA98 : dout <= 12'h131;
		12'hA99 : dout <= 12'h12F;
		12'hA9A : dout <= 12'h12D;
		12'hA9B : dout <= 12'h12C;
		12'hA9C : dout <= 12'h12A;
		12'hA9D : dout <= 12'h129;
		12'hA9E : dout <= 12'h127;
		12'hA9F : dout <= 12'h125;
		12'hAA0 : dout <= 12'h124;
		12'hAA1 : dout <= 12'h122;
		12'hAA2 : dout <= 12'h121;
		12'hAA3 : dout <= 12'h11F;
		12'hAA4 : dout <= 12'h11D;
		12'hAA5 : dout <= 12'h11C;
		12'hAA6 : dout <= 12'h11A;
		12'hAA7 : dout <= 12'h119;
		12'hAA8 : dout <= 12'h117;
		12'hAA9 : dout <= 12'h115;
		12'hAAA : dout <= 12'h114;
		12'hAAB : dout <= 12'h112;
		12'hAAC : dout <= 12'h111;
		12'hAAD : dout <= 12'h10F;
		12'hAAE : dout <= 12'h10E;
		12'hAAF : dout <= 12'h10C;
		12'hAB0 : dout <= 12'h10A;
		12'hAB1 : dout <= 12'h109;
		12'hAB2 : dout <= 12'h107;
		12'hAB3 : dout <= 12'h106;
		12'hAB4 : dout <= 12'h104;
		12'hAB5 : dout <= 12'h103;
		12'hAB6 : dout <= 12'h101;
		12'hAB7 : dout <= 12'h100;
		12'hAB8 : dout <= 12'h0FE;
		12'hAB9 : dout <= 12'h0FD;
		12'hABA : dout <= 12'h0FB;
		12'hABB : dout <= 12'h0FA;
		12'hABC : dout <= 12'h0F8;
		12'hABD : dout <= 12'h0F7;
		12'hABE : dout <= 12'h0F5;
		12'hABF : dout <= 12'h0F4;
		12'hAC0 : dout <= 12'h0F2;
		12'hAC1 : dout <= 12'h0F1;
		12'hAC2 : dout <= 12'h0EF;
		12'hAC3 : dout <= 12'h0EE;
		12'hAC4 : dout <= 12'h0EC;
		12'hAC5 : dout <= 12'h0EB;
		12'hAC6 : dout <= 12'h0E9;
		12'hAC7 : dout <= 12'h0E8;
		12'hAC8 : dout <= 12'h0E7;
		12'hAC9 : dout <= 12'h0E5;
		12'hACA : dout <= 12'h0E4;
		12'hACB : dout <= 12'h0E2;
		12'hACC : dout <= 12'h0E1;
		12'hACD : dout <= 12'h0DF;
		12'hACE : dout <= 12'h0DE;
		12'hACF : dout <= 12'h0DC;
		12'hAD0 : dout <= 12'h0DB;
		12'hAD1 : dout <= 12'h0DA;
		12'hAD2 : dout <= 12'h0D8;
		12'hAD3 : dout <= 12'h0D7;
		12'hAD4 : dout <= 12'h0D5;
		12'hAD5 : dout <= 12'h0D4;
		12'hAD6 : dout <= 12'h0D3;
		12'hAD7 : dout <= 12'h0D1;
		12'hAD8 : dout <= 12'h0D0;
		12'hAD9 : dout <= 12'h0CF;
		12'hADA : dout <= 12'h0CD;
		12'hADB : dout <= 12'h0CC;
		12'hADC : dout <= 12'h0CA;
		12'hADD : dout <= 12'h0C9;
		12'hADE : dout <= 12'h0C8;
		12'hADF : dout <= 12'h0C6;
		12'hAE0 : dout <= 12'h0C5;
		12'hAE1 : dout <= 12'h0C4;
		12'hAE2 : dout <= 12'h0C2;
		12'hAE3 : dout <= 12'h0C1;
		12'hAE4 : dout <= 12'h0C0;
		12'hAE5 : dout <= 12'h0BE;
		12'hAE6 : dout <= 12'h0BD;
		12'hAE7 : dout <= 12'h0BC;
		12'hAE8 : dout <= 12'h0BA;
		12'hAE9 : dout <= 12'h0B9;
		12'hAEA : dout <= 12'h0B8;
		12'hAEB : dout <= 12'h0B7;
		12'hAEC : dout <= 12'h0B5;
		12'hAED : dout <= 12'h0B4;
		12'hAEE : dout <= 12'h0B3;
		12'hAEF : dout <= 12'h0B1;
		12'hAF0 : dout <= 12'h0B0;
		12'hAF1 : dout <= 12'h0AF;
		12'hAF2 : dout <= 12'h0AE;
		12'hAF3 : dout <= 12'h0AC;
		12'hAF4 : dout <= 12'h0AB;
		12'hAF5 : dout <= 12'h0AA;
		12'hAF6 : dout <= 12'h0A9;
		12'hAF7 : dout <= 12'h0A7;
		12'hAF8 : dout <= 12'h0A6;
		12'hAF9 : dout <= 12'h0A5;
		12'hAFA : dout <= 12'h0A4;
		12'hAFB : dout <= 12'h0A2;
		12'hAFC : dout <= 12'h0A1;
		12'hAFD : dout <= 12'h0A0;
		12'hAFE : dout <= 12'h09F;
		12'hAFF : dout <= 12'h09E;
		12'hB00 : dout <= 12'h09C;
		12'hB01 : dout <= 12'h09B;
		12'hB02 : dout <= 12'h09A;
		12'hB03 : dout <= 12'h099;
		12'hB04 : dout <= 12'h098;
		12'hB05 : dout <= 12'h096;
		12'hB06 : dout <= 12'h095;
		12'hB07 : dout <= 12'h094;
		12'hB08 : dout <= 12'h093;
		12'hB09 : dout <= 12'h092;
		12'hB0A : dout <= 12'h091;
		12'hB0B : dout <= 12'h08F;
		12'hB0C : dout <= 12'h08E;
		12'hB0D : dout <= 12'h08D;
		12'hB0E : dout <= 12'h08C;
		12'hB0F : dout <= 12'h08B;
		12'hB10 : dout <= 12'h08A;
		12'hB11 : dout <= 12'h089;
		12'hB12 : dout <= 12'h087;
		12'hB13 : dout <= 12'h086;
		12'hB14 : dout <= 12'h085;
		12'hB15 : dout <= 12'h084;
		12'hB16 : dout <= 12'h083;
		12'hB17 : dout <= 12'h082;
		12'hB18 : dout <= 12'h081;
		12'hB19 : dout <= 12'h080;
		12'hB1A : dout <= 12'h07F;
		12'hB1B : dout <= 12'h07E;
		12'hB1C : dout <= 12'h07C;
		12'hB1D : dout <= 12'h07B;
		12'hB1E : dout <= 12'h07A;
		12'hB1F : dout <= 12'h079;
		12'hB20 : dout <= 12'h078;
		12'hB21 : dout <= 12'h077;
		12'hB22 : dout <= 12'h076;
		12'hB23 : dout <= 12'h075;
		12'hB24 : dout <= 12'h074;
		12'hB25 : dout <= 12'h073;
		12'hB26 : dout <= 12'h072;
		12'hB27 : dout <= 12'h071;
		12'hB28 : dout <= 12'h070;
		12'hB29 : dout <= 12'h06F;
		12'hB2A : dout <= 12'h06E;
		12'hB2B : dout <= 12'h06D;
		12'hB2C : dout <= 12'h06C;
		12'hB2D : dout <= 12'h06B;
		12'hB2E : dout <= 12'h06A;
		12'hB2F : dout <= 12'h069;
		12'hB30 : dout <= 12'h068;
		12'hB31 : dout <= 12'h067;
		12'hB32 : dout <= 12'h066;
		12'hB33 : dout <= 12'h065;
		12'hB34 : dout <= 12'h064;
		12'hB35 : dout <= 12'h063;
		12'hB36 : dout <= 12'h062;
		12'hB37 : dout <= 12'h061;
		12'hB38 : dout <= 12'h060;
		12'hB39 : dout <= 12'h05F;
		12'hB3A : dout <= 12'h05E;
		12'hB3B : dout <= 12'h05D;
		12'hB3C : dout <= 12'h05C;
		12'hB3D : dout <= 12'h05B;
		12'hB3E : dout <= 12'h05A;
		12'hB3F : dout <= 12'h05A;
		12'hB40 : dout <= 12'h059;
		12'hB41 : dout <= 12'h058;
		12'hB42 : dout <= 12'h057;
		12'hB43 : dout <= 12'h056;
		12'hB44 : dout <= 12'h055;
		12'hB45 : dout <= 12'h054;
		12'hB46 : dout <= 12'h053;
		12'hB47 : dout <= 12'h052;
		12'hB48 : dout <= 12'h051;
		12'hB49 : dout <= 12'h051;
		12'hB4A : dout <= 12'h050;
		12'hB4B : dout <= 12'h04F;
		12'hB4C : dout <= 12'h04E;
		12'hB4D : dout <= 12'h04D;
		12'hB4E : dout <= 12'h04C;
		12'hB4F : dout <= 12'h04B;
		12'hB50 : dout <= 12'h04B;
		12'hB51 : dout <= 12'h04A;
		12'hB52 : dout <= 12'h049;
		12'hB53 : dout <= 12'h048;
		12'hB54 : dout <= 12'h047;
		12'hB55 : dout <= 12'h047;
		12'hB56 : dout <= 12'h046;
		12'hB57 : dout <= 12'h045;
		12'hB58 : dout <= 12'h044;
		12'hB59 : dout <= 12'h043;
		12'hB5A : dout <= 12'h043;
		12'hB5B : dout <= 12'h042;
		12'hB5C : dout <= 12'h041;
		12'hB5D : dout <= 12'h040;
		12'hB5E : dout <= 12'h03F;
		12'hB5F : dout <= 12'h03F;
		12'hB60 : dout <= 12'h03E;
		12'hB61 : dout <= 12'h03D;
		12'hB62 : dout <= 12'h03C;
		12'hB63 : dout <= 12'h03C;
		12'hB64 : dout <= 12'h03B;
		12'hB65 : dout <= 12'h03A;
		12'hB66 : dout <= 12'h039;
		12'hB67 : dout <= 12'h039;
		12'hB68 : dout <= 12'h038;
		12'hB69 : dout <= 12'h037;
		12'hB6A : dout <= 12'h036;
		12'hB6B : dout <= 12'h036;
		12'hB6C : dout <= 12'h035;
		12'hB6D : dout <= 12'h034;
		12'hB6E : dout <= 12'h034;
		12'hB6F : dout <= 12'h033;
		12'hB70 : dout <= 12'h032;
		12'hB71 : dout <= 12'h032;
		12'hB72 : dout <= 12'h031;
		12'hB73 : dout <= 12'h030;
		12'hB74 : dout <= 12'h030;
		12'hB75 : dout <= 12'h02F;
		12'hB76 : dout <= 12'h02E;
		12'hB77 : dout <= 12'h02E;
		12'hB78 : dout <= 12'h02D;
		12'hB79 : dout <= 12'h02C;
		12'hB7A : dout <= 12'h02C;
		12'hB7B : dout <= 12'h02B;
		12'hB7C : dout <= 12'h02A;
		12'hB7D : dout <= 12'h02A;
		12'hB7E : dout <= 12'h029;
		12'hB7F : dout <= 12'h028;
		12'hB80 : dout <= 12'h028;
		12'hB81 : dout <= 12'h027;
		12'hB82 : dout <= 12'h027;
		12'hB83 : dout <= 12'h026;
		12'hB84 : dout <= 12'h025;
		12'hB85 : dout <= 12'h025;
		12'hB86 : dout <= 12'h024;
		12'hB87 : dout <= 12'h024;
		12'hB88 : dout <= 12'h023;
		12'hB89 : dout <= 12'h023;
		12'hB8A : dout <= 12'h022;
		12'hB8B : dout <= 12'h021;
		12'hB8C : dout <= 12'h021;
		12'hB8D : dout <= 12'h020;
		12'hB8E : dout <= 12'h020;
		12'hB8F : dout <= 12'h01F;
		12'hB90 : dout <= 12'h01F;
		12'hB91 : dout <= 12'h01E;
		12'hB92 : dout <= 12'h01E;
		12'hB93 : dout <= 12'h01D;
		12'hB94 : dout <= 12'h01D;
		12'hB95 : dout <= 12'h01C;
		12'hB96 : dout <= 12'h01C;
		12'hB97 : dout <= 12'h01B;
		12'hB98 : dout <= 12'h01A;
		12'hB99 : dout <= 12'h01A;
		12'hB9A : dout <= 12'h01A;
		12'hB9B : dout <= 12'h019;
		12'hB9C : dout <= 12'h019;
		12'hB9D : dout <= 12'h018;
		12'hB9E : dout <= 12'h018;
		12'hB9F : dout <= 12'h017;
		12'hBA0 : dout <= 12'h017;
		12'hBA1 : dout <= 12'h016;
		12'hBA2 : dout <= 12'h016;
		12'hBA3 : dout <= 12'h015;
		12'hBA4 : dout <= 12'h015;
		12'hBA5 : dout <= 12'h014;
		12'hBA6 : dout <= 12'h014;
		12'hBA7 : dout <= 12'h014;
		12'hBA8 : dout <= 12'h013;
		12'hBA9 : dout <= 12'h013;
		12'hBAA : dout <= 12'h012;
		12'hBAB : dout <= 12'h012;
		12'hBAC : dout <= 12'h011;
		12'hBAD : dout <= 12'h011;
		12'hBAE : dout <= 12'h011;
		12'hBAF : dout <= 12'h010;
		12'hBB0 : dout <= 12'h010;
		12'hBB1 : dout <= 12'h010;
		12'hBB2 : dout <= 12'h00F;
		12'hBB3 : dout <= 12'h00F;
		12'hBB4 : dout <= 12'h00E;
		12'hBB5 : dout <= 12'h00E;
		12'hBB6 : dout <= 12'h00E;
		12'hBB7 : dout <= 12'h00D;
		12'hBB8 : dout <= 12'h00D;
		12'hBB9 : dout <= 12'h00D;
		12'hBBA : dout <= 12'h00C;
		12'hBBB : dout <= 12'h00C;
		12'hBBC : dout <= 12'h00C;
		12'hBBD : dout <= 12'h00B;
		12'hBBE : dout <= 12'h00B;
		12'hBBF : dout <= 12'h00B;
		12'hBC0 : dout <= 12'h00A;
		12'hBC1 : dout <= 12'h00A;
		12'hBC2 : dout <= 12'h00A;
		12'hBC3 : dout <= 12'h009;
		12'hBC4 : dout <= 12'h009;
		12'hBC5 : dout <= 12'h009;
		12'hBC6 : dout <= 12'h009;
		12'hBC7 : dout <= 12'h008;
		12'hBC8 : dout <= 12'h008;
		12'hBC9 : dout <= 12'h008;
		12'hBCA : dout <= 12'h008;
		12'hBCB : dout <= 12'h007;
		12'hBCC : dout <= 12'h007;
		12'hBCD : dout <= 12'h007;
		12'hBCE : dout <= 12'h007;
		12'hBCF : dout <= 12'h006;
		12'hBD0 : dout <= 12'h006;
		12'hBD1 : dout <= 12'h006;
		12'hBD2 : dout <= 12'h006;
		12'hBD3 : dout <= 12'h005;
		12'hBD4 : dout <= 12'h005;
		12'hBD5 : dout <= 12'h005;
		12'hBD6 : dout <= 12'h005;
		12'hBD7 : dout <= 12'h005;
		12'hBD8 : dout <= 12'h004;
		12'hBD9 : dout <= 12'h004;
		12'hBDA : dout <= 12'h004;
		12'hBDB : dout <= 12'h004;
		12'hBDC : dout <= 12'h004;
		12'hBDD : dout <= 12'h003;
		12'hBDE : dout <= 12'h003;
		12'hBDF : dout <= 12'h003;
		12'hBE0 : dout <= 12'h003;
		12'hBE1 : dout <= 12'h003;
		12'hBE2 : dout <= 12'h003;
		12'hBE3 : dout <= 12'h003;
		12'hBE4 : dout <= 12'h002;
		12'hBE5 : dout <= 12'h002;
		12'hBE6 : dout <= 12'h002;
		12'hBE7 : dout <= 12'h002;
		12'hBE8 : dout <= 12'h002;
		12'hBE9 : dout <= 12'h002;
		12'hBEA : dout <= 12'h002;
		12'hBEB : dout <= 12'h002;
		12'hBEC : dout <= 12'h001;
		12'hBED : dout <= 12'h001;
		12'hBEE : dout <= 12'h001;
		12'hBEF : dout <= 12'h001;
		12'hBF0 : dout <= 12'h001;
		12'hBF1 : dout <= 12'h001;
		12'hBF2 : dout <= 12'h001;
		12'hBF3 : dout <= 12'h001;
		12'hBF4 : dout <= 12'h001;
		12'hBF5 : dout <= 12'h001;
		12'hBF6 : dout <= 12'h001;
		12'hBF7 : dout <= 12'h001;
		12'hBF8 : dout <= 12'h001;
		12'hBF9 : dout <= 12'h001;
		12'hBFA : dout <= 12'h001;
		12'hBFB : dout <= 12'h001;
		12'hBFC : dout <= 12'h001;
		12'hBFD : dout <= 12'h001;
		12'hBFE : dout <= 12'h001;
		12'hBFF : dout <= 12'h001;
		12'hC00 : dout <= 12'h000;
		12'hC01 : dout <= 12'h001;
		12'hC02 : dout <= 12'h001;
		12'hC03 : dout <= 12'h001;
		12'hC04 : dout <= 12'h001;
		12'hC05 : dout <= 12'h001;
		12'hC06 : dout <= 12'h001;
		12'hC07 : dout <= 12'h001;
		12'hC08 : dout <= 12'h001;
		12'hC09 : dout <= 12'h001;
		12'hC0A : dout <= 12'h001;
		12'hC0B : dout <= 12'h001;
		12'hC0C : dout <= 12'h001;
		12'hC0D : dout <= 12'h001;
		12'hC0E : dout <= 12'h001;
		12'hC0F : dout <= 12'h001;
		12'hC10 : dout <= 12'h001;
		12'hC11 : dout <= 12'h001;
		12'hC12 : dout <= 12'h001;
		12'hC13 : dout <= 12'h001;
		12'hC14 : dout <= 12'h001;
		12'hC15 : dout <= 12'h002;
		12'hC16 : dout <= 12'h002;
		12'hC17 : dout <= 12'h002;
		12'hC18 : dout <= 12'h002;
		12'hC19 : dout <= 12'h002;
		12'hC1A : dout <= 12'h002;
		12'hC1B : dout <= 12'h002;
		12'hC1C : dout <= 12'h002;
		12'hC1D : dout <= 12'h003;
		12'hC1E : dout <= 12'h003;
		12'hC1F : dout <= 12'h003;
		12'hC20 : dout <= 12'h003;
		12'hC21 : dout <= 12'h003;
		12'hC22 : dout <= 12'h003;
		12'hC23 : dout <= 12'h003;
		12'hC24 : dout <= 12'h004;
		12'hC25 : dout <= 12'h004;
		12'hC26 : dout <= 12'h004;
		12'hC27 : dout <= 12'h004;
		12'hC28 : dout <= 12'h004;
		12'hC29 : dout <= 12'h005;
		12'hC2A : dout <= 12'h005;
		12'hC2B : dout <= 12'h005;
		12'hC2C : dout <= 12'h005;
		12'hC2D : dout <= 12'h005;
		12'hC2E : dout <= 12'h006;
		12'hC2F : dout <= 12'h006;
		12'hC30 : dout <= 12'h006;
		12'hC31 : dout <= 12'h006;
		12'hC32 : dout <= 12'h007;
		12'hC33 : dout <= 12'h007;
		12'hC34 : dout <= 12'h007;
		12'hC35 : dout <= 12'h007;
		12'hC36 : dout <= 12'h008;
		12'hC37 : dout <= 12'h008;
		12'hC38 : dout <= 12'h008;
		12'hC39 : dout <= 12'h008;
		12'hC3A : dout <= 12'h009;
		12'hC3B : dout <= 12'h009;
		12'hC3C : dout <= 12'h009;
		12'hC3D : dout <= 12'h009;
		12'hC3E : dout <= 12'h00A;
		12'hC3F : dout <= 12'h00A;
		12'hC40 : dout <= 12'h00A;
		12'hC41 : dout <= 12'h00B;
		12'hC42 : dout <= 12'h00B;
		12'hC43 : dout <= 12'h00B;
		12'hC44 : dout <= 12'h00C;
		12'hC45 : dout <= 12'h00C;
		12'hC46 : dout <= 12'h00C;
		12'hC47 : dout <= 12'h00D;
		12'hC48 : dout <= 12'h00D;
		12'hC49 : dout <= 12'h00D;
		12'hC4A : dout <= 12'h00E;
		12'hC4B : dout <= 12'h00E;
		12'hC4C : dout <= 12'h00E;
		12'hC4D : dout <= 12'h00F;
		12'hC4E : dout <= 12'h00F;
		12'hC4F : dout <= 12'h010;
		12'hC50 : dout <= 12'h010;
		12'hC51 : dout <= 12'h010;
		12'hC52 : dout <= 12'h011;
		12'hC53 : dout <= 12'h011;
		12'hC54 : dout <= 12'h011;
		12'hC55 : dout <= 12'h012;
		12'hC56 : dout <= 12'h012;
		12'hC57 : dout <= 12'h013;
		12'hC58 : dout <= 12'h013;
		12'hC59 : dout <= 12'h014;
		12'hC5A : dout <= 12'h014;
		12'hC5B : dout <= 12'h014;
		12'hC5C : dout <= 12'h015;
		12'hC5D : dout <= 12'h015;
		12'hC5E : dout <= 12'h016;
		12'hC5F : dout <= 12'h016;
		12'hC60 : dout <= 12'h017;
		12'hC61 : dout <= 12'h017;
		12'hC62 : dout <= 12'h018;
		12'hC63 : dout <= 12'h018;
		12'hC64 : dout <= 12'h019;
		12'hC65 : dout <= 12'h019;
		12'hC66 : dout <= 12'h01A;
		12'hC67 : dout <= 12'h01A;
		12'hC68 : dout <= 12'h01A;
		12'hC69 : dout <= 12'h01B;
		12'hC6A : dout <= 12'h01C;
		12'hC6B : dout <= 12'h01C;
		12'hC6C : dout <= 12'h01D;
		12'hC6D : dout <= 12'h01D;
		12'hC6E : dout <= 12'h01E;
		12'hC6F : dout <= 12'h01E;
		12'hC70 : dout <= 12'h01F;
		12'hC71 : dout <= 12'h01F;
		12'hC72 : dout <= 12'h020;
		12'hC73 : dout <= 12'h020;
		12'hC74 : dout <= 12'h021;
		12'hC75 : dout <= 12'h021;
		12'hC76 : dout <= 12'h022;
		12'hC77 : dout <= 12'h023;
		12'hC78 : dout <= 12'h023;
		12'hC79 : dout <= 12'h024;
		12'hC7A : dout <= 12'h024;
		12'hC7B : dout <= 12'h025;
		12'hC7C : dout <= 12'h025;
		12'hC7D : dout <= 12'h026;
		12'hC7E : dout <= 12'h027;
		12'hC7F : dout <= 12'h027;
		12'hC80 : dout <= 12'h028;
		12'hC81 : dout <= 12'h028;
		12'hC82 : dout <= 12'h029;
		12'hC83 : dout <= 12'h02A;
		12'hC84 : dout <= 12'h02A;
		12'hC85 : dout <= 12'h02B;
		12'hC86 : dout <= 12'h02C;
		12'hC87 : dout <= 12'h02C;
		12'hC88 : dout <= 12'h02D;
		12'hC89 : dout <= 12'h02E;
		12'hC8A : dout <= 12'h02E;
		12'hC8B : dout <= 12'h02F;
		12'hC8C : dout <= 12'h030;
		12'hC8D : dout <= 12'h030;
		12'hC8E : dout <= 12'h031;
		12'hC8F : dout <= 12'h032;
		12'hC90 : dout <= 12'h032;
		12'hC91 : dout <= 12'h033;
		12'hC92 : dout <= 12'h034;
		12'hC93 : dout <= 12'h034;
		12'hC94 : dout <= 12'h035;
		12'hC95 : dout <= 12'h036;
		12'hC96 : dout <= 12'h036;
		12'hC97 : dout <= 12'h037;
		12'hC98 : dout <= 12'h038;
		12'hC99 : dout <= 12'h039;
		12'hC9A : dout <= 12'h039;
		12'hC9B : dout <= 12'h03A;
		12'hC9C : dout <= 12'h03B;
		12'hC9D : dout <= 12'h03C;
		12'hC9E : dout <= 12'h03C;
		12'hC9F : dout <= 12'h03D;
		12'hCA0 : dout <= 12'h03E;
		12'hCA1 : dout <= 12'h03F;
		12'hCA2 : dout <= 12'h03F;
		12'hCA3 : dout <= 12'h040;
		12'hCA4 : dout <= 12'h041;
		12'hCA5 : dout <= 12'h042;
		12'hCA6 : dout <= 12'h043;
		12'hCA7 : dout <= 12'h043;
		12'hCA8 : dout <= 12'h044;
		12'hCA9 : dout <= 12'h045;
		12'hCAA : dout <= 12'h046;
		12'hCAB : dout <= 12'h047;
		12'hCAC : dout <= 12'h047;
		12'hCAD : dout <= 12'h048;
		12'hCAE : dout <= 12'h049;
		12'hCAF : dout <= 12'h04A;
		12'hCB0 : dout <= 12'h04B;
		12'hCB1 : dout <= 12'h04B;
		12'hCB2 : dout <= 12'h04C;
		12'hCB3 : dout <= 12'h04D;
		12'hCB4 : dout <= 12'h04E;
		12'hCB5 : dout <= 12'h04F;
		12'hCB6 : dout <= 12'h050;
		12'hCB7 : dout <= 12'h051;
		12'hCB8 : dout <= 12'h051;
		12'hCB9 : dout <= 12'h052;
		12'hCBA : dout <= 12'h053;
		12'hCBB : dout <= 12'h054;
		12'hCBC : dout <= 12'h055;
		12'hCBD : dout <= 12'h056;
		12'hCBE : dout <= 12'h057;
		12'hCBF : dout <= 12'h058;
		12'hCC0 : dout <= 12'h059;
		12'hCC1 : dout <= 12'h05A;
		12'hCC2 : dout <= 12'h05A;
		12'hCC3 : dout <= 12'h05B;
		12'hCC4 : dout <= 12'h05C;
		12'hCC5 : dout <= 12'h05D;
		12'hCC6 : dout <= 12'h05E;
		12'hCC7 : dout <= 12'h05F;
		12'hCC8 : dout <= 12'h060;
		12'hCC9 : dout <= 12'h061;
		12'hCCA : dout <= 12'h062;
		12'hCCB : dout <= 12'h063;
		12'hCCC : dout <= 12'h064;
		12'hCCD : dout <= 12'h065;
		12'hCCE : dout <= 12'h066;
		12'hCCF : dout <= 12'h067;
		12'hCD0 : dout <= 12'h068;
		12'hCD1 : dout <= 12'h069;
		12'hCD2 : dout <= 12'h06A;
		12'hCD3 : dout <= 12'h06B;
		12'hCD4 : dout <= 12'h06C;
		12'hCD5 : dout <= 12'h06D;
		12'hCD6 : dout <= 12'h06E;
		12'hCD7 : dout <= 12'h06F;
		12'hCD8 : dout <= 12'h070;
		12'hCD9 : dout <= 12'h071;
		12'hCDA : dout <= 12'h072;
		12'hCDB : dout <= 12'h073;
		12'hCDC : dout <= 12'h074;
		12'hCDD : dout <= 12'h075;
		12'hCDE : dout <= 12'h076;
		12'hCDF : dout <= 12'h077;
		12'hCE0 : dout <= 12'h078;
		12'hCE1 : dout <= 12'h079;
		12'hCE2 : dout <= 12'h07A;
		12'hCE3 : dout <= 12'h07B;
		12'hCE4 : dout <= 12'h07C;
		12'hCE5 : dout <= 12'h07E;
		12'hCE6 : dout <= 12'h07F;
		12'hCE7 : dout <= 12'h080;
		12'hCE8 : dout <= 12'h081;
		12'hCE9 : dout <= 12'h082;
		12'hCEA : dout <= 12'h083;
		12'hCEB : dout <= 12'h084;
		12'hCEC : dout <= 12'h085;
		12'hCED : dout <= 12'h086;
		12'hCEE : dout <= 12'h087;
		12'hCEF : dout <= 12'h089;
		12'hCF0 : dout <= 12'h08A;
		12'hCF1 : dout <= 12'h08B;
		12'hCF2 : dout <= 12'h08C;
		12'hCF3 : dout <= 12'h08D;
		12'hCF4 : dout <= 12'h08E;
		12'hCF5 : dout <= 12'h08F;
		12'hCF6 : dout <= 12'h091;
		12'hCF7 : dout <= 12'h092;
		12'hCF8 : dout <= 12'h093;
		12'hCF9 : dout <= 12'h094;
		12'hCFA : dout <= 12'h095;
		12'hCFB : dout <= 12'h096;
		12'hCFC : dout <= 12'h098;
		12'hCFD : dout <= 12'h099;
		12'hCFE : dout <= 12'h09A;
		12'hCFF : dout <= 12'h09B;
		12'hD00 : dout <= 12'h09C;
		12'hD01 : dout <= 12'h09E;
		12'hD02 : dout <= 12'h09F;
		12'hD03 : dout <= 12'h0A0;
		12'hD04 : dout <= 12'h0A1;
		12'hD05 : dout <= 12'h0A2;
		12'hD06 : dout <= 12'h0A4;
		12'hD07 : dout <= 12'h0A5;
		12'hD08 : dout <= 12'h0A6;
		12'hD09 : dout <= 12'h0A7;
		12'hD0A : dout <= 12'h0A9;
		12'hD0B : dout <= 12'h0AA;
		12'hD0C : dout <= 12'h0AB;
		12'hD0D : dout <= 12'h0AC;
		12'hD0E : dout <= 12'h0AE;
		12'hD0F : dout <= 12'h0AF;
		12'hD10 : dout <= 12'h0B0;
		12'hD11 : dout <= 12'h0B1;
		12'hD12 : dout <= 12'h0B3;
		12'hD13 : dout <= 12'h0B4;
		12'hD14 : dout <= 12'h0B5;
		12'hD15 : dout <= 12'h0B7;
		12'hD16 : dout <= 12'h0B8;
		12'hD17 : dout <= 12'h0B9;
		12'hD18 : dout <= 12'h0BA;
		12'hD19 : dout <= 12'h0BC;
		12'hD1A : dout <= 12'h0BD;
		12'hD1B : dout <= 12'h0BE;
		12'hD1C : dout <= 12'h0C0;
		12'hD1D : dout <= 12'h0C1;
		12'hD1E : dout <= 12'h0C2;
		12'hD1F : dout <= 12'h0C4;
		12'hD20 : dout <= 12'h0C5;
		12'hD21 : dout <= 12'h0C6;
		12'hD22 : dout <= 12'h0C8;
		12'hD23 : dout <= 12'h0C9;
		12'hD24 : dout <= 12'h0CA;
		12'hD25 : dout <= 12'h0CC;
		12'hD26 : dout <= 12'h0CD;
		12'hD27 : dout <= 12'h0CF;
		12'hD28 : dout <= 12'h0D0;
		12'hD29 : dout <= 12'h0D1;
		12'hD2A : dout <= 12'h0D3;
		12'hD2B : dout <= 12'h0D4;
		12'hD2C : dout <= 12'h0D5;
		12'hD2D : dout <= 12'h0D7;
		12'hD2E : dout <= 12'h0D8;
		12'hD2F : dout <= 12'h0DA;
		12'hD30 : dout <= 12'h0DB;
		12'hD31 : dout <= 12'h0DC;
		12'hD32 : dout <= 12'h0DE;
		12'hD33 : dout <= 12'h0DF;
		12'hD34 : dout <= 12'h0E1;
		12'hD35 : dout <= 12'h0E2;
		12'hD36 : dout <= 12'h0E4;
		12'hD37 : dout <= 12'h0E5;
		12'hD38 : dout <= 12'h0E7;
		12'hD39 : dout <= 12'h0E8;
		12'hD3A : dout <= 12'h0E9;
		12'hD3B : dout <= 12'h0EB;
		12'hD3C : dout <= 12'h0EC;
		12'hD3D : dout <= 12'h0EE;
		12'hD3E : dout <= 12'h0EF;
		12'hD3F : dout <= 12'h0F1;
		12'hD40 : dout <= 12'h0F2;
		12'hD41 : dout <= 12'h0F4;
		12'hD42 : dout <= 12'h0F5;
		12'hD43 : dout <= 12'h0F7;
		12'hD44 : dout <= 12'h0F8;
		12'hD45 : dout <= 12'h0FA;
		12'hD46 : dout <= 12'h0FB;
		12'hD47 : dout <= 12'h0FD;
		12'hD48 : dout <= 12'h0FE;
		12'hD49 : dout <= 12'h100;
		12'hD4A : dout <= 12'h101;
		12'hD4B : dout <= 12'h103;
		12'hD4C : dout <= 12'h104;
		12'hD4D : dout <= 12'h106;
		12'hD4E : dout <= 12'h107;
		12'hD4F : dout <= 12'h109;
		12'hD50 : dout <= 12'h10A;
		12'hD51 : dout <= 12'h10C;
		12'hD52 : dout <= 12'h10E;
		12'hD53 : dout <= 12'h10F;
		12'hD54 : dout <= 12'h111;
		12'hD55 : dout <= 12'h112;
		12'hD56 : dout <= 12'h114;
		12'hD57 : dout <= 12'h115;
		12'hD58 : dout <= 12'h117;
		12'hD59 : dout <= 12'h119;
		12'hD5A : dout <= 12'h11A;
		12'hD5B : dout <= 12'h11C;
		12'hD5C : dout <= 12'h11D;
		12'hD5D : dout <= 12'h11F;
		12'hD5E : dout <= 12'h121;
		12'hD5F : dout <= 12'h122;
		12'hD60 : dout <= 12'h124;
		12'hD61 : dout <= 12'h125;
		12'hD62 : dout <= 12'h127;
		12'hD63 : dout <= 12'h129;
		12'hD64 : dout <= 12'h12A;
		12'hD65 : dout <= 12'h12C;
		12'hD66 : dout <= 12'h12D;
		12'hD67 : dout <= 12'h12F;
		12'hD68 : dout <= 12'h131;
		12'hD69 : dout <= 12'h132;
		12'hD6A : dout <= 12'h134;
		12'hD6B : dout <= 12'h136;
		12'hD6C : dout <= 12'h137;
		12'hD6D : dout <= 12'h139;
		12'hD6E : dout <= 12'h13B;
		12'hD6F : dout <= 12'h13C;
		12'hD70 : dout <= 12'h13E;
		12'hD71 : dout <= 12'h140;
		12'hD72 : dout <= 12'h141;
		12'hD73 : dout <= 12'h143;
		12'hD74 : dout <= 12'h145;
		12'hD75 : dout <= 12'h147;
		12'hD76 : dout <= 12'h148;
		12'hD77 : dout <= 12'h14A;
		12'hD78 : dout <= 12'h14C;
		12'hD79 : dout <= 12'h14D;
		12'hD7A : dout <= 12'h14F;
		12'hD7B : dout <= 12'h151;
		12'hD7C : dout <= 12'h153;
		12'hD7D : dout <= 12'h154;
		12'hD7E : dout <= 12'h156;
		12'hD7F : dout <= 12'h158;
		12'hD80 : dout <= 12'h159;
		12'hD81 : dout <= 12'h15B;
		12'hD82 : dout <= 12'h15D;
		12'hD83 : dout <= 12'h15F;
		12'hD84 : dout <= 12'h160;
		12'hD85 : dout <= 12'h162;
		12'hD86 : dout <= 12'h164;
		12'hD87 : dout <= 12'h166;
		12'hD88 : dout <= 12'h168;
		12'hD89 : dout <= 12'h169;
		12'hD8A : dout <= 12'h16B;
		12'hD8B : dout <= 12'h16D;
		12'hD8C : dout <= 12'h16F;
		12'hD8D : dout <= 12'h170;
		12'hD8E : dout <= 12'h172;
		12'hD8F : dout <= 12'h174;
		12'hD90 : dout <= 12'h176;
		12'hD91 : dout <= 12'h178;
		12'hD92 : dout <= 12'h17A;
		12'hD93 : dout <= 12'h17B;
		12'hD94 : dout <= 12'h17D;
		12'hD95 : dout <= 12'h17F;
		12'hD96 : dout <= 12'h181;
		12'hD97 : dout <= 12'h183;
		12'hD98 : dout <= 12'h184;
		12'hD99 : dout <= 12'h186;
		12'hD9A : dout <= 12'h188;
		12'hD9B : dout <= 12'h18A;
		12'hD9C : dout <= 12'h18C;
		12'hD9D : dout <= 12'h18E;
		12'hD9E : dout <= 12'h190;
		12'hD9F : dout <= 12'h191;
		12'hDA0 : dout <= 12'h193;
		12'hDA1 : dout <= 12'h195;
		12'hDA2 : dout <= 12'h197;
		12'hDA3 : dout <= 12'h199;
		12'hDA4 : dout <= 12'h19B;
		12'hDA5 : dout <= 12'h19D;
		12'hDA6 : dout <= 12'h19F;
		12'hDA7 : dout <= 12'h1A1;
		12'hDA8 : dout <= 12'h1A2;
		12'hDA9 : dout <= 12'h1A4;
		12'hDAA : dout <= 12'h1A6;
		12'hDAB : dout <= 12'h1A8;
		12'hDAC : dout <= 12'h1AA;
		12'hDAD : dout <= 12'h1AC;
		12'hDAE : dout <= 12'h1AE;
		12'hDAF : dout <= 12'h1B0;
		12'hDB0 : dout <= 12'h1B2;
		12'hDB1 : dout <= 12'h1B4;
		12'hDB2 : dout <= 12'h1B6;
		12'hDB3 : dout <= 12'h1B8;
		12'hDB4 : dout <= 12'h1BA;
		12'hDB5 : dout <= 12'h1BB;
		12'hDB6 : dout <= 12'h1BD;
		12'hDB7 : dout <= 12'h1BF;
		12'hDB8 : dout <= 12'h1C1;
		12'hDB9 : dout <= 12'h1C3;
		12'hDBA : dout <= 12'h1C5;
		12'hDBB : dout <= 12'h1C7;
		12'hDBC : dout <= 12'h1C9;
		12'hDBD : dout <= 12'h1CB;
		12'hDBE : dout <= 12'h1CD;
		12'hDBF : dout <= 12'h1CF;
		12'hDC0 : dout <= 12'h1D1;
		12'hDC1 : dout <= 12'h1D3;
		12'hDC2 : dout <= 12'h1D5;
		12'hDC3 : dout <= 12'h1D7;
		12'hDC4 : dout <= 12'h1D9;
		12'hDC5 : dout <= 12'h1DB;
		12'hDC6 : dout <= 12'h1DD;
		12'hDC7 : dout <= 12'h1DF;
		12'hDC8 : dout <= 12'h1E1;
		12'hDC9 : dout <= 12'h1E3;
		12'hDCA : dout <= 12'h1E5;
		12'hDCB : dout <= 12'h1E7;
		12'hDCC : dout <= 12'h1E9;
		12'hDCD : dout <= 12'h1EB;
		12'hDCE : dout <= 12'h1ED;
		12'hDCF : dout <= 12'h1EF;
		12'hDD0 : dout <= 12'h1F1;
		12'hDD1 : dout <= 12'h1F4;
		12'hDD2 : dout <= 12'h1F6;
		12'hDD3 : dout <= 12'h1F8;
		12'hDD4 : dout <= 12'h1FA;
		12'hDD5 : dout <= 12'h1FC;
		12'hDD6 : dout <= 12'h1FE;
		12'hDD7 : dout <= 12'h200;
		12'hDD8 : dout <= 12'h202;
		12'hDD9 : dout <= 12'h204;
		12'hDDA : dout <= 12'h206;
		12'hDDB : dout <= 12'h208;
		12'hDDC : dout <= 12'h20A;
		12'hDDD : dout <= 12'h20C;
		12'hDDE : dout <= 12'h20F;
		12'hDDF : dout <= 12'h211;
		12'hDE0 : dout <= 12'h213;
		12'hDE1 : dout <= 12'h215;
		12'hDE2 : dout <= 12'h217;
		12'hDE3 : dout <= 12'h219;
		12'hDE4 : dout <= 12'h21B;
		12'hDE5 : dout <= 12'h21D;
		12'hDE6 : dout <= 12'h21F;
		12'hDE7 : dout <= 12'h222;
		12'hDE8 : dout <= 12'h224;
		12'hDE9 : dout <= 12'h226;
		12'hDEA : dout <= 12'h228;
		12'hDEB : dout <= 12'h22A;
		12'hDEC : dout <= 12'h22C;
		12'hDED : dout <= 12'h22E;
		12'hDEE : dout <= 12'h231;
		12'hDEF : dout <= 12'h233;
		12'hDF0 : dout <= 12'h235;
		12'hDF1 : dout <= 12'h237;
		12'hDF2 : dout <= 12'h239;
		12'hDF3 : dout <= 12'h23B;
		12'hDF4 : dout <= 12'h23E;
		12'hDF5 : dout <= 12'h240;
		12'hDF6 : dout <= 12'h242;
		12'hDF7 : dout <= 12'h244;
		12'hDF8 : dout <= 12'h246;
		12'hDF9 : dout <= 12'h249;
		12'hDFA : dout <= 12'h24B;
		12'hDFB : dout <= 12'h24D;
		12'hDFC : dout <= 12'h24F;
		12'hDFD : dout <= 12'h251;
		12'hDFE : dout <= 12'h254;
		12'hDFF : dout <= 12'h256;
		12'hE00 : dout <= 12'h258;
		12'hE01 : dout <= 12'h25A;
		12'hE02 : dout <= 12'h25C;
		12'hE03 : dout <= 12'h25F;
		12'hE04 : dout <= 12'h261;
		12'hE05 : dout <= 12'h263;
		12'hE06 : dout <= 12'h265;
		12'hE07 : dout <= 12'h268;
		12'hE08 : dout <= 12'h26A;
		12'hE09 : dout <= 12'h26C;
		12'hE0A : dout <= 12'h26E;
		12'hE0B : dout <= 12'h271;
		12'hE0C : dout <= 12'h273;
		12'hE0D : dout <= 12'h275;
		12'hE0E : dout <= 12'h277;
		12'hE0F : dout <= 12'h27A;
		12'hE10 : dout <= 12'h27C;
		12'hE11 : dout <= 12'h27E;
		12'hE12 : dout <= 12'h281;
		12'hE13 : dout <= 12'h283;
		12'hE14 : dout <= 12'h285;
		12'hE15 : dout <= 12'h287;
		12'hE16 : dout <= 12'h28A;
		12'hE17 : dout <= 12'h28C;
		12'hE18 : dout <= 12'h28E;
		12'hE19 : dout <= 12'h291;
		12'hE1A : dout <= 12'h293;
		12'hE1B : dout <= 12'h295;
		12'hE1C : dout <= 12'h298;
		12'hE1D : dout <= 12'h29A;
		12'hE1E : dout <= 12'h29C;
		12'hE1F : dout <= 12'h29E;
		12'hE20 : dout <= 12'h2A1;
		12'hE21 : dout <= 12'h2A3;
		12'hE22 : dout <= 12'h2A5;
		12'hE23 : dout <= 12'h2A8;
		12'hE24 : dout <= 12'h2AA;
		12'hE25 : dout <= 12'h2AC;
		12'hE26 : dout <= 12'h2AF;
		12'hE27 : dout <= 12'h2B1;
		12'hE28 : dout <= 12'h2B4;
		12'hE29 : dout <= 12'h2B6;
		12'hE2A : dout <= 12'h2B8;
		12'hE2B : dout <= 12'h2BB;
		12'hE2C : dout <= 12'h2BD;
		12'hE2D : dout <= 12'h2BF;
		12'hE2E : dout <= 12'h2C2;
		12'hE2F : dout <= 12'h2C4;
		12'hE30 : dout <= 12'h2C6;
		12'hE31 : dout <= 12'h2C9;
		12'hE32 : dout <= 12'h2CB;
		12'hE33 : dout <= 12'h2CE;
		12'hE34 : dout <= 12'h2D0;
		12'hE35 : dout <= 12'h2D2;
		12'hE36 : dout <= 12'h2D5;
		12'hE37 : dout <= 12'h2D7;
		12'hE38 : dout <= 12'h2DA;
		12'hE39 : dout <= 12'h2DC;
		12'hE3A : dout <= 12'h2DE;
		12'hE3B : dout <= 12'h2E1;
		12'hE3C : dout <= 12'h2E3;
		12'hE3D : dout <= 12'h2E6;
		12'hE3E : dout <= 12'h2E8;
		12'hE3F : dout <= 12'h2EA;
		12'hE40 : dout <= 12'h2ED;
		12'hE41 : dout <= 12'h2EF;
		12'hE42 : dout <= 12'h2F2;
		12'hE43 : dout <= 12'h2F4;
		12'hE44 : dout <= 12'h2F7;
		12'hE45 : dout <= 12'h2F9;
		12'hE46 : dout <= 12'h2FC;
		12'hE47 : dout <= 12'h2FE;
		12'hE48 : dout <= 12'h300;
		12'hE49 : dout <= 12'h303;
		12'hE4A : dout <= 12'h305;
		12'hE4B : dout <= 12'h308;
		12'hE4C : dout <= 12'h30A;
		12'hE4D : dout <= 12'h30D;
		12'hE4E : dout <= 12'h30F;
		12'hE4F : dout <= 12'h312;
		12'hE50 : dout <= 12'h314;
		12'hE51 : dout <= 12'h317;
		12'hE52 : dout <= 12'h319;
		12'hE53 : dout <= 12'h31C;
		12'hE54 : dout <= 12'h31E;
		12'hE55 : dout <= 12'h321;
		12'hE56 : dout <= 12'h323;
		12'hE57 : dout <= 12'h326;
		12'hE58 : dout <= 12'h328;
		12'hE59 : dout <= 12'h32B;
		12'hE5A : dout <= 12'h32D;
		12'hE5B : dout <= 12'h330;
		12'hE5C : dout <= 12'h332;
		12'hE5D : dout <= 12'h335;
		12'hE5E : dout <= 12'h337;
		12'hE5F : dout <= 12'h33A;
		12'hE60 : dout <= 12'h33C;
		12'hE61 : dout <= 12'h33F;
		12'hE62 : dout <= 12'h341;
		12'hE63 : dout <= 12'h344;
		12'hE64 : dout <= 12'h346;
		12'hE65 : dout <= 12'h349;
		12'hE66 : dout <= 12'h34B;
		12'hE67 : dout <= 12'h34E;
		12'hE68 : dout <= 12'h350;
		12'hE69 : dout <= 12'h353;
		12'hE6A : dout <= 12'h355;
		12'hE6B : dout <= 12'h358;
		12'hE6C : dout <= 12'h35B;
		12'hE6D : dout <= 12'h35D;
		12'hE6E : dout <= 12'h360;
		12'hE6F : dout <= 12'h362;
		12'hE70 : dout <= 12'h365;
		12'hE71 : dout <= 12'h367;
		12'hE72 : dout <= 12'h36A;
		12'hE73 : dout <= 12'h36D;
		12'hE74 : dout <= 12'h36F;
		12'hE75 : dout <= 12'h372;
		12'hE76 : dout <= 12'h374;
		12'hE77 : dout <= 12'h377;
		12'hE78 : dout <= 12'h379;
		12'hE79 : dout <= 12'h37C;
		12'hE7A : dout <= 12'h37F;
		12'hE7B : dout <= 12'h381;
		12'hE7C : dout <= 12'h384;
		12'hE7D : dout <= 12'h386;
		12'hE7E : dout <= 12'h389;
		12'hE7F : dout <= 12'h38C;
		12'hE80 : dout <= 12'h38E;
		12'hE81 : dout <= 12'h391;
		12'hE82 : dout <= 12'h393;
		12'hE83 : dout <= 12'h396;
		12'hE84 : dout <= 12'h399;
		12'hE85 : dout <= 12'h39B;
		12'hE86 : dout <= 12'h39E;
		12'hE87 : dout <= 12'h3A1;
		12'hE88 : dout <= 12'h3A3;
		12'hE89 : dout <= 12'h3A6;
		12'hE8A : dout <= 12'h3A8;
		12'hE8B : dout <= 12'h3AB;
		12'hE8C : dout <= 12'h3AE;
		12'hE8D : dout <= 12'h3B0;
		12'hE8E : dout <= 12'h3B3;
		12'hE8F : dout <= 12'h3B6;
		12'hE90 : dout <= 12'h3B8;
		12'hE91 : dout <= 12'h3BB;
		12'hE92 : dout <= 12'h3BE;
		12'hE93 : dout <= 12'h3C0;
		12'hE94 : dout <= 12'h3C3;
		12'hE95 : dout <= 12'h3C6;
		12'hE96 : dout <= 12'h3C8;
		12'hE97 : dout <= 12'h3CB;
		12'hE98 : dout <= 12'h3CE;
		12'hE99 : dout <= 12'h3D0;
		12'hE9A : dout <= 12'h3D3;
		12'hE9B : dout <= 12'h3D6;
		12'hE9C : dout <= 12'h3D8;
		12'hE9D : dout <= 12'h3DB;
		12'hE9E : dout <= 12'h3DE;
		12'hE9F : dout <= 12'h3E0;
		12'hEA0 : dout <= 12'h3E3;
		12'hEA1 : dout <= 12'h3E6;
		12'hEA2 : dout <= 12'h3E9;
		12'hEA3 : dout <= 12'h3EB;
		12'hEA4 : dout <= 12'h3EE;
		12'hEA5 : dout <= 12'h3F1;
		12'hEA6 : dout <= 12'h3F3;
		12'hEA7 : dout <= 12'h3F6;
		12'hEA8 : dout <= 12'h3F9;
		12'hEA9 : dout <= 12'h3FB;
		12'hEAA : dout <= 12'h3FE;
		12'hEAB : dout <= 12'h401;
		12'hEAC : dout <= 12'h404;
		12'hEAD : dout <= 12'h406;
		12'hEAE : dout <= 12'h409;
		12'hEAF : dout <= 12'h40C;
		12'hEB0 : dout <= 12'h40F;
		12'hEB1 : dout <= 12'h411;
		12'hEB2 : dout <= 12'h414;
		12'hEB3 : dout <= 12'h417;
		12'hEB4 : dout <= 12'h419;
		12'hEB5 : dout <= 12'h41C;
		12'hEB6 : dout <= 12'h41F;
		12'hEB7 : dout <= 12'h422;
		12'hEB8 : dout <= 12'h424;
		12'hEB9 : dout <= 12'h427;
		12'hEBA : dout <= 12'h42A;
		12'hEBB : dout <= 12'h42D;
		12'hEBC : dout <= 12'h42F;
		12'hEBD : dout <= 12'h432;
		12'hEBE : dout <= 12'h435;
		12'hEBF : dout <= 12'h438;
		12'hEC0 : dout <= 12'h43B;
		12'hEC1 : dout <= 12'h43D;
		12'hEC2 : dout <= 12'h440;
		12'hEC3 : dout <= 12'h443;
		12'hEC4 : dout <= 12'h446;
		12'hEC5 : dout <= 12'h448;
		12'hEC6 : dout <= 12'h44B;
		12'hEC7 : dout <= 12'h44E;
		12'hEC8 : dout <= 12'h451;
		12'hEC9 : dout <= 12'h454;
		12'hECA : dout <= 12'h456;
		12'hECB : dout <= 12'h459;
		12'hECC : dout <= 12'h45C;
		12'hECD : dout <= 12'h45F;
		12'hECE : dout <= 12'h462;
		12'hECF : dout <= 12'h464;
		12'hED0 : dout <= 12'h467;
		12'hED1 : dout <= 12'h46A;
		12'hED2 : dout <= 12'h46D;
		12'hED3 : dout <= 12'h470;
		12'hED4 : dout <= 12'h472;
		12'hED5 : dout <= 12'h475;
		12'hED6 : dout <= 12'h478;
		12'hED7 : dout <= 12'h47B;
		12'hED8 : dout <= 12'h47E;
		12'hED9 : dout <= 12'h480;
		12'hEDA : dout <= 12'h483;
		12'hEDB : dout <= 12'h486;
		12'hEDC : dout <= 12'h489;
		12'hEDD : dout <= 12'h48C;
		12'hEDE : dout <= 12'h48F;
		12'hEDF : dout <= 12'h491;
		12'hEE0 : dout <= 12'h494;
		12'hEE1 : dout <= 12'h497;
		12'hEE2 : dout <= 12'h49A;
		12'hEE3 : dout <= 12'h49D;
		12'hEE4 : dout <= 12'h4A0;
		12'hEE5 : dout <= 12'h4A3;
		12'hEE6 : dout <= 12'h4A5;
		12'hEE7 : dout <= 12'h4A8;
		12'hEE8 : dout <= 12'h4AB;
		12'hEE9 : dout <= 12'h4AE;
		12'hEEA : dout <= 12'h4B1;
		12'hEEB : dout <= 12'h4B4;
		12'hEEC : dout <= 12'h4B7;
		12'hEED : dout <= 12'h4B9;
		12'hEEE : dout <= 12'h4BC;
		12'hEEF : dout <= 12'h4BF;
		12'hEF0 : dout <= 12'h4C2;
		12'hEF1 : dout <= 12'h4C5;
		12'hEF2 : dout <= 12'h4C8;
		12'hEF3 : dout <= 12'h4CB;
		12'hEF4 : dout <= 12'h4CD;
		12'hEF5 : dout <= 12'h4D0;
		12'hEF6 : dout <= 12'h4D3;
		12'hEF7 : dout <= 12'h4D6;
		12'hEF8 : dout <= 12'h4D9;
		12'hEF9 : dout <= 12'h4DC;
		12'hEFA : dout <= 12'h4DF;
		12'hEFB : dout <= 12'h4E2;
		12'hEFC : dout <= 12'h4E5;
		12'hEFD : dout <= 12'h4E7;
		12'hEFE : dout <= 12'h4EA;
		12'hEFF : dout <= 12'h4ED;
		12'hF00 : dout <= 12'h4F0;
		12'hF01 : dout <= 12'h4F3;
		12'hF02 : dout <= 12'h4F6;
		12'hF03 : dout <= 12'h4F9;
		12'hF04 : dout <= 12'h4FC;
		12'hF05 : dout <= 12'h4FF;
		12'hF06 : dout <= 12'h502;
		12'hF07 : dout <= 12'h504;
		12'hF08 : dout <= 12'h507;
		12'hF09 : dout <= 12'h50A;
		12'hF0A : dout <= 12'h50D;
		12'hF0B : dout <= 12'h510;
		12'hF0C : dout <= 12'h513;
		12'hF0D : dout <= 12'h516;
		12'hF0E : dout <= 12'h519;
		12'hF0F : dout <= 12'h51C;
		12'hF10 : dout <= 12'h51F;
		12'hF11 : dout <= 12'h522;
		12'hF12 : dout <= 12'h525;
		12'hF13 : dout <= 12'h528;
		12'hF14 : dout <= 12'h52B;
		12'hF15 : dout <= 12'h52D;
		12'hF16 : dout <= 12'h530;
		12'hF17 : dout <= 12'h533;
		12'hF18 : dout <= 12'h536;
		12'hF19 : dout <= 12'h539;
		12'hF1A : dout <= 12'h53C;
		12'hF1B : dout <= 12'h53F;
		12'hF1C : dout <= 12'h542;
		12'hF1D : dout <= 12'h545;
		12'hF1E : dout <= 12'h548;
		12'hF1F : dout <= 12'h54B;
		12'hF20 : dout <= 12'h54E;
		12'hF21 : dout <= 12'h551;
		12'hF22 : dout <= 12'h554;
		12'hF23 : dout <= 12'h557;
		12'hF24 : dout <= 12'h55A;
		12'hF25 : dout <= 12'h55D;
		12'hF26 : dout <= 12'h560;
		12'hF27 : dout <= 12'h563;
		12'hF28 : dout <= 12'h566;
		12'hF29 : dout <= 12'h569;
		12'hF2A : dout <= 12'h56C;
		12'hF2B : dout <= 12'h56F;
		12'hF2C : dout <= 12'h571;
		12'hF2D : dout <= 12'h574;
		12'hF2E : dout <= 12'h577;
		12'hF2F : dout <= 12'h57A;
		12'hF30 : dout <= 12'h57D;
		12'hF31 : dout <= 12'h580;
		12'hF32 : dout <= 12'h583;
		12'hF33 : dout <= 12'h586;
		12'hF34 : dout <= 12'h589;
		12'hF35 : dout <= 12'h58C;
		12'hF36 : dout <= 12'h58F;
		12'hF37 : dout <= 12'h592;
		12'hF38 : dout <= 12'h595;
		12'hF39 : dout <= 12'h598;
		12'hF3A : dout <= 12'h59B;
		12'hF3B : dout <= 12'h59E;
		12'hF3C : dout <= 12'h5A1;
		12'hF3D : dout <= 12'h5A4;
		12'hF3E : dout <= 12'h5A7;
		12'hF3F : dout <= 12'h5AA;
		12'hF40 : dout <= 12'h5AD;
		12'hF41 : dout <= 12'h5B0;
		12'hF42 : dout <= 12'h5B3;
		12'hF43 : dout <= 12'h5B6;
		12'hF44 : dout <= 12'h5B9;
		12'hF45 : dout <= 12'h5BC;
		12'hF46 : dout <= 12'h5BF;
		12'hF47 : dout <= 12'h5C2;
		12'hF48 : dout <= 12'h5C5;
		12'hF49 : dout <= 12'h5C8;
		12'hF4A : dout <= 12'h5CB;
		12'hF4B : dout <= 12'h5CE;
		12'hF4C : dout <= 12'h5D1;
		12'hF4D : dout <= 12'h5D4;
		12'hF4E : dout <= 12'h5D7;
		12'hF4F : dout <= 12'h5DB;
		12'hF50 : dout <= 12'h5DE;
		12'hF51 : dout <= 12'h5E1;
		12'hF52 : dout <= 12'h5E4;
		12'hF53 : dout <= 12'h5E7;
		12'hF54 : dout <= 12'h5EA;
		12'hF55 : dout <= 12'h5ED;
		12'hF56 : dout <= 12'h5F0;
		12'hF57 : dout <= 12'h5F3;
		12'hF58 : dout <= 12'h5F6;
		12'hF59 : dout <= 12'h5F9;
		12'hF5A : dout <= 12'h5FC;
		12'hF5B : dout <= 12'h5FF;
		12'hF5C : dout <= 12'h602;
		12'hF5D : dout <= 12'h605;
		12'hF5E : dout <= 12'h608;
		12'hF5F : dout <= 12'h60B;
		12'hF60 : dout <= 12'h60E;
		12'hF61 : dout <= 12'h611;
		12'hF62 : dout <= 12'h614;
		12'hF63 : dout <= 12'h617;
		12'hF64 : dout <= 12'h61A;
		12'hF65 : dout <= 12'h61D;
		12'hF66 : dout <= 12'h620;
		12'hF67 : dout <= 12'h623;
		12'hF68 : dout <= 12'h627;
		12'hF69 : dout <= 12'h62A;
		12'hF6A : dout <= 12'h62D;
		12'hF6B : dout <= 12'h630;
		12'hF6C : dout <= 12'h633;
		12'hF6D : dout <= 12'h636;
		12'hF6E : dout <= 12'h639;
		12'hF6F : dout <= 12'h63C;
		12'hF70 : dout <= 12'h63F;
		12'hF71 : dout <= 12'h642;
		12'hF72 : dout <= 12'h645;
		12'hF73 : dout <= 12'h648;
		12'hF74 : dout <= 12'h64B;
		12'hF75 : dout <= 12'h64E;
		12'hF76 : dout <= 12'h651;
		12'hF77 : dout <= 12'h654;
		12'hF78 : dout <= 12'h658;
		12'hF79 : dout <= 12'h65B;
		12'hF7A : dout <= 12'h65E;
		12'hF7B : dout <= 12'h661;
		12'hF7C : dout <= 12'h664;
		12'hF7D : dout <= 12'h667;
		12'hF7E : dout <= 12'h66A;
		12'hF7F : dout <= 12'h66D;
		12'hF80 : dout <= 12'h670;
		12'hF81 : dout <= 12'h673;
		12'hF82 : dout <= 12'h676;
		12'hF83 : dout <= 12'h679;
		12'hF84 : dout <= 12'h67C;
		12'hF85 : dout <= 12'h680;
		12'hF86 : dout <= 12'h683;
		12'hF87 : dout <= 12'h686;
		12'hF88 : dout <= 12'h689;
		12'hF89 : dout <= 12'h68C;
		12'hF8A : dout <= 12'h68F;
		12'hF8B : dout <= 12'h692;
		12'hF8C : dout <= 12'h695;
		12'hF8D : dout <= 12'h698;
		12'hF8E : dout <= 12'h69B;
		12'hF8F : dout <= 12'h69E;
		12'hF90 : dout <= 12'h6A2;
		12'hF91 : dout <= 12'h6A5;
		12'hF92 : dout <= 12'h6A8;
		12'hF93 : dout <= 12'h6AB;
		12'hF94 : dout <= 12'h6AE;
		12'hF95 : dout <= 12'h6B1;
		12'hF96 : dout <= 12'h6B4;
		12'hF97 : dout <= 12'h6B7;
		12'hF98 : dout <= 12'h6BA;
		12'hF99 : dout <= 12'h6BD;
		12'hF9A : dout <= 12'h6C1;
		12'hF9B : dout <= 12'h6C4;
		12'hF9C : dout <= 12'h6C7;
		12'hF9D : dout <= 12'h6CA;
		12'hF9E : dout <= 12'h6CD;
		12'hF9F : dout <= 12'h6D0;
		12'hFA0 : dout <= 12'h6D3;
		12'hFA1 : dout <= 12'h6D6;
		12'hFA2 : dout <= 12'h6D9;
		12'hFA3 : dout <= 12'h6DC;
		12'hFA4 : dout <= 12'h6E0;
		12'hFA5 : dout <= 12'h6E3;
		12'hFA6 : dout <= 12'h6E6;
		12'hFA7 : dout <= 12'h6E9;
		12'hFA8 : dout <= 12'h6EC;
		12'hFA9 : dout <= 12'h6EF;
		12'hFAA : dout <= 12'h6F2;
		12'hFAB : dout <= 12'h6F5;
		12'hFAC : dout <= 12'h6F8;
		12'hFAD : dout <= 12'h6FC;
		12'hFAE : dout <= 12'h6FF;
		12'hFAF : dout <= 12'h702;
		12'hFB0 : dout <= 12'h705;
		12'hFB1 : dout <= 12'h708;
		12'hFB2 : dout <= 12'h70B;
		12'hFB3 : dout <= 12'h70E;
		12'hFB4 : dout <= 12'h711;
		12'hFB5 : dout <= 12'h715;
		12'hFB6 : dout <= 12'h718;
		12'hFB7 : dout <= 12'h71B;
		12'hFB8 : dout <= 12'h71E;
		12'hFB9 : dout <= 12'h721;
		12'hFBA : dout <= 12'h724;
		12'hFBB : dout <= 12'h727;
		12'hFBC : dout <= 12'h72A;
		12'hFBD : dout <= 12'h72D;
		12'hFBE : dout <= 12'h731;
		12'hFBF : dout <= 12'h734;
		12'hFC0 : dout <= 12'h737;
		12'hFC1 : dout <= 12'h73A;
		12'hFC2 : dout <= 12'h73D;
		12'hFC3 : dout <= 12'h740;
		12'hFC4 : dout <= 12'h743;
		12'hFC5 : dout <= 12'h746;
		12'hFC6 : dout <= 12'h74A;
		12'hFC7 : dout <= 12'h74D;
		12'hFC8 : dout <= 12'h750;
		12'hFC9 : dout <= 12'h753;
		12'hFCA : dout <= 12'h756;
		12'hFCB : dout <= 12'h759;
		12'hFCC : dout <= 12'h75C;
		12'hFCD : dout <= 12'h760;
		12'hFCE : dout <= 12'h763;
		12'hFCF : dout <= 12'h766;
		12'hFD0 : dout <= 12'h769;
		12'hFD1 : dout <= 12'h76C;
		12'hFD2 : dout <= 12'h76F;
		12'hFD3 : dout <= 12'h772;
		12'hFD4 : dout <= 12'h775;
		12'hFD5 : dout <= 12'h779;
		12'hFD6 : dout <= 12'h77C;
		12'hFD7 : dout <= 12'h77F;
		12'hFD8 : dout <= 12'h782;
		12'hFD9 : dout <= 12'h785;
		12'hFDA : dout <= 12'h788;
		12'hFDB : dout <= 12'h78B;
		12'hFDC : dout <= 12'h78F;
		12'hFDD : dout <= 12'h792;
		12'hFDE : dout <= 12'h795;
		12'hFDF : dout <= 12'h798;
		12'hFE0 : dout <= 12'h79B;
		12'hFE1 : dout <= 12'h79E;
		12'hFE2 : dout <= 12'h7A1;
		12'hFE3 : dout <= 12'h7A4;
		12'hFE4 : dout <= 12'h7A8;
		12'hFE5 : dout <= 12'h7AB;
		12'hFE6 : dout <= 12'h7AE;
		12'hFE7 : dout <= 12'h7B1;
		12'hFE8 : dout <= 12'h7B4;
		12'hFE9 : dout <= 12'h7B7;
		12'hFEA : dout <= 12'h7BA;
		12'hFEB : dout <= 12'h7BE;
		12'hFEC : dout <= 12'h7C1;
		12'hFED : dout <= 12'h7C4;
		12'hFEE : dout <= 12'h7C7;
		12'hFEF : dout <= 12'h7CA;
		12'hFF0 : dout <= 12'h7CD;
		12'hFF1 : dout <= 12'h7D0;
		12'hFF2 : dout <= 12'h7D4;
		12'hFF3 : dout <= 12'h7D7;
		12'hFF4 : dout <= 12'h7DA;
		12'hFF5 : dout <= 12'h7DD;
		12'hFF6 : dout <= 12'h7E0;
		12'hFF7 : dout <= 12'h7E3;
		12'hFF8 : dout <= 12'h7E6;
		12'hFF9 : dout <= 12'h7EA;
		12'hFFA : dout <= 12'h7ED;
		12'hFFB : dout <= 12'h7F0;
		12'hFFC : dout <= 12'h7F3;
		12'hFFD : dout <= 12'h7F6;
		12'hFFE : dout <= 12'h7F9;
		12'hFFF : dout <= 12'h7FC;
		endcase
end	

endmodule