module usin_rom
(
	input			clk		,
	input			rst 	,
	input	[11:0]	addr	,

	output	[11:0]	dout
);
		
	always@ (posedge clk, negedge rst) begin
		if (!rst)
			dout_r <= 0;
		else
			case (addr)
			12'h000 : dout_r <= 12'h800;
			12'h001 : dout_r <= 12'h803;
			12'h002 : dout_r <= 12'h806;
			12'h003 : dout_r <= 12'h809;
			12'h004 : dout_r <= 12'h80C;
			12'h005 : dout_r <= 12'h80F;
			12'h006 : dout_r <= 12'h812;
			12'h007 : dout_r <= 12'h815;
			12'h008 : dout_r <= 12'h819;
			12'h009 : dout_r <= 12'h81C;
			12'h00A : dout_r <= 12'h81F;
			12'h00B : dout_r <= 12'h822;
			12'h00C : dout_r <= 12'h825;
			12'h00D : dout_r <= 12'h828;
			12'h00E : dout_r <= 12'h82B;
			12'h00F : dout_r <= 12'h82F;
			12'h010 : dout_r <= 12'h832;
			12'h011 : dout_r <= 12'h835;
			12'h012 : dout_r <= 12'h838;
			12'h013 : dout_r <= 12'h83B;
			12'h014 : dout_r <= 12'h83E;
			12'h015 : dout_r <= 12'h841;
			12'h016 : dout_r <= 12'h845;
			12'h017 : dout_r <= 12'h848;
			12'h018 : dout_r <= 12'h84B;
			12'h019 : dout_r <= 12'h84E;
			12'h01A : dout_r <= 12'h851;
			12'h01B : dout_r <= 12'h854;
			12'h01C : dout_r <= 12'h857;
			12'h01D : dout_r <= 12'h85B;
			12'h01E : dout_r <= 12'h85E;
			12'h01F : dout_r <= 12'h861;
			12'h020 : dout_r <= 12'h864;
			12'h021 : dout_r <= 12'h867;
			12'h022 : dout_r <= 12'h86A;
			12'h023 : dout_r <= 12'h86D;
			12'h024 : dout_r <= 12'h870;
			12'h025 : dout_r <= 12'h874;
			12'h026 : dout_r <= 12'h877;
			12'h027 : dout_r <= 12'h87A;
			12'h028 : dout_r <= 12'h87D;
			12'h029 : dout_r <= 12'h880;
			12'h02A : dout_r <= 12'h883;
			12'h02B : dout_r <= 12'h886;
			12'h02C : dout_r <= 12'h88A;
			12'h02D : dout_r <= 12'h88D;
			12'h02E : dout_r <= 12'h890;
			12'h02F : dout_r <= 12'h893;
			12'h030 : dout_r <= 12'h896;
			12'h031 : dout_r <= 12'h899;
			12'h032 : dout_r <= 12'h89C;
			12'h033 : dout_r <= 12'h89F;
			12'h034 : dout_r <= 12'h8A3;
			12'h035 : dout_r <= 12'h8A6;
			12'h036 : dout_r <= 12'h8A9;
			12'h037 : dout_r <= 12'h8AC;
			12'h038 : dout_r <= 12'h8AF;
			12'h039 : dout_r <= 12'h8B2;
			12'h03A : dout_r <= 12'h8B5;
			12'h03B : dout_r <= 12'h8B9;
			12'h03C : dout_r <= 12'h8BC;
			12'h03D : dout_r <= 12'h8BF;
			12'h03E : dout_r <= 12'h8C2;
			12'h03F : dout_r <= 12'h8C5;
			12'h040 : dout_r <= 12'h8C8;
			12'h041 : dout_r <= 12'h8CB;
			12'h042 : dout_r <= 12'h8CE;
			12'h043 : dout_r <= 12'h8D2;
			12'h044 : dout_r <= 12'h8D5;
			12'h045 : dout_r <= 12'h8D8;
			12'h046 : dout_r <= 12'h8DB;
			12'h047 : dout_r <= 12'h8DE;
			12'h048 : dout_r <= 12'h8E1;
			12'h049 : dout_r <= 12'h8E4;
			12'h04A : dout_r <= 12'h8E7;
			12'h04B : dout_r <= 12'h8EA;
			12'h04C : dout_r <= 12'h8EE;
			12'h04D : dout_r <= 12'h8F1;
			12'h04E : dout_r <= 12'h8F4;
			12'h04F : dout_r <= 12'h8F7;
			12'h050 : dout_r <= 12'h8FA;
			12'h051 : dout_r <= 12'h8FD;
			12'h052 : dout_r <= 12'h900;
			12'h053 : dout_r <= 12'h903;
			12'h054 : dout_r <= 12'h907;
			12'h055 : dout_r <= 12'h90A;
			12'h056 : dout_r <= 12'h90D;
			12'h057 : dout_r <= 12'h910;
			12'h058 : dout_r <= 12'h913;
			12'h059 : dout_r <= 12'h916;
			12'h05A : dout_r <= 12'h919;
			12'h05B : dout_r <= 12'h91C;
			12'h05C : dout_r <= 12'h91F;
			12'h05D : dout_r <= 12'h923;
			12'h05E : dout_r <= 12'h926;
			12'h05F : dout_r <= 12'h929;
			12'h060 : dout_r <= 12'h92C;
			12'h061 : dout_r <= 12'h92F;
			12'h062 : dout_r <= 12'h932;
			12'h063 : dout_r <= 12'h935;
			12'h064 : dout_r <= 12'h938;
			12'h065 : dout_r <= 12'h93B;
			12'h066 : dout_r <= 12'h93E;
			12'h067 : dout_r <= 12'h942;
			12'h068 : dout_r <= 12'h945;
			12'h069 : dout_r <= 12'h948;
			12'h06A : dout_r <= 12'h94B;
			12'h06B : dout_r <= 12'h94E;
			12'h06C : dout_r <= 12'h951;
			12'h06D : dout_r <= 12'h954;
			12'h06E : dout_r <= 12'h957;
			12'h06F : dout_r <= 12'h95A;
			12'h070 : dout_r <= 12'h95D;
			12'h071 : dout_r <= 12'h961;
			12'h072 : dout_r <= 12'h964;
			12'h073 : dout_r <= 12'h967;
			12'h074 : dout_r <= 12'h96A;
			12'h075 : dout_r <= 12'h96D;
			12'h076 : dout_r <= 12'h970;
			12'h077 : dout_r <= 12'h973;
			12'h078 : dout_r <= 12'h976;
			12'h079 : dout_r <= 12'h979;
			12'h07A : dout_r <= 12'h97C;
			12'h07B : dout_r <= 12'h97F;
			12'h07C : dout_r <= 12'h983;
			12'h07D : dout_r <= 12'h986;
			12'h07E : dout_r <= 12'h989;
			12'h07F : dout_r <= 12'h98C;
			12'h080 : dout_r <= 12'h98F;
			12'h081 : dout_r <= 12'h992;
			12'h082 : dout_r <= 12'h995;
			12'h083 : dout_r <= 12'h998;
			12'h084 : dout_r <= 12'h99B;
			12'h085 : dout_r <= 12'h99E;
			12'h086 : dout_r <= 12'h9A1;
			12'h087 : dout_r <= 12'h9A4;
			12'h088 : dout_r <= 12'h9A7;
			12'h089 : dout_r <= 12'h9AB;
			12'h08A : dout_r <= 12'h9AE;
			12'h08B : dout_r <= 12'h9B1;
			12'h08C : dout_r <= 12'h9B4;
			12'h08D : dout_r <= 12'h9B7;
			12'h08E : dout_r <= 12'h9BA;
			12'h08F : dout_r <= 12'h9BD;
			12'h090 : dout_r <= 12'h9C0;
			12'h091 : dout_r <= 12'h9C3;
			12'h092 : dout_r <= 12'h9C6;
			12'h093 : dout_r <= 12'h9C9;
			12'h094 : dout_r <= 12'h9CC;
			12'h095 : dout_r <= 12'h9CF;
			12'h096 : dout_r <= 12'h9D2;
			12'h097 : dout_r <= 12'h9D5;
			12'h098 : dout_r <= 12'h9D8;
			12'h099 : dout_r <= 12'h9DC;
			12'h09A : dout_r <= 12'h9DF;
			12'h09B : dout_r <= 12'h9E2;
			12'h09C : dout_r <= 12'h9E5;
			12'h09D : dout_r <= 12'h9E8;
			12'h09E : dout_r <= 12'h9EB;
			12'h09F : dout_r <= 12'h9EE;
			12'h0A0 : dout_r <= 12'h9F1;
			12'h0A1 : dout_r <= 12'h9F4;
			12'h0A2 : dout_r <= 12'h9F7;
			12'h0A3 : dout_r <= 12'h9FA;
			12'h0A4 : dout_r <= 12'h9FD;
			12'h0A5 : dout_r <= 12'hA00;
			12'h0A6 : dout_r <= 12'hA03;
			12'h0A7 : dout_r <= 12'hA06;
			12'h0A8 : dout_r <= 12'hA09;
			12'h0A9 : dout_r <= 12'hA0C;
			12'h0AA : dout_r <= 12'hA0F;
			12'h0AB : dout_r <= 12'hA12;
			12'h0AC : dout_r <= 12'hA15;
			12'h0AD : dout_r <= 12'hA18;
			12'h0AE : dout_r <= 12'hA1B;
			12'h0AF : dout_r <= 12'hA1E;
			12'h0B0 : dout_r <= 12'hA21;
			12'h0B1 : dout_r <= 12'hA24;
			12'h0B2 : dout_r <= 12'hA28;
			12'h0B3 : dout_r <= 12'hA2B;
			12'h0B4 : dout_r <= 12'hA2E;
			12'h0B5 : dout_r <= 12'hA31;
			12'h0B6 : dout_r <= 12'hA34;
			12'h0B7 : dout_r <= 12'hA37;
			12'h0B8 : dout_r <= 12'hA3A;
			12'h0B9 : dout_r <= 12'hA3D;
			12'h0BA : dout_r <= 12'hA40;
			12'h0BB : dout_r <= 12'hA43;
			12'h0BC : dout_r <= 12'hA46;
			12'h0BD : dout_r <= 12'hA49;
			12'h0BE : dout_r <= 12'hA4C;
			12'h0BF : dout_r <= 12'hA4F;
			12'h0C0 : dout_r <= 12'hA52;
			12'h0C1 : dout_r <= 12'hA55;
			12'h0C2 : dout_r <= 12'hA58;
			12'h0C3 : dout_r <= 12'hA5B;
			12'h0C4 : dout_r <= 12'hA5E;
			12'h0C5 : dout_r <= 12'hA61;
			12'h0C6 : dout_r <= 12'hA64;
			12'h0C7 : dout_r <= 12'hA67;
			12'h0C8 : dout_r <= 12'hA6A;
			12'h0C9 : dout_r <= 12'hA6D;
			12'h0CA : dout_r <= 12'hA70;
			12'h0CB : dout_r <= 12'hA73;
			12'h0CC : dout_r <= 12'hA76;
			12'h0CD : dout_r <= 12'hA79;
			12'h0CE : dout_r <= 12'hA7C;
			12'h0CF : dout_r <= 12'hA7F;
			12'h0D0 : dout_r <= 12'hA82;
			12'h0D1 : dout_r <= 12'hA85;
			12'h0D2 : dout_r <= 12'hA88;
			12'h0D3 : dout_r <= 12'hA8B;
			12'h0D4 : dout_r <= 12'hA8E;
			12'h0D5 : dout_r <= 12'hA90;
			12'h0D6 : dout_r <= 12'hA93;
			12'h0D7 : dout_r <= 12'hA96;
			12'h0D8 : dout_r <= 12'hA99;
			12'h0D9 : dout_r <= 12'hA9C;
			12'h0DA : dout_r <= 12'hA9F;
			12'h0DB : dout_r <= 12'hAA2;
			12'h0DC : dout_r <= 12'hAA5;
			12'h0DD : dout_r <= 12'hAA8;
			12'h0DE : dout_r <= 12'hAAB;
			12'h0DF : dout_r <= 12'hAAE;
			12'h0E0 : dout_r <= 12'hAB1;
			12'h0E1 : dout_r <= 12'hAB4;
			12'h0E2 : dout_r <= 12'hAB7;
			12'h0E3 : dout_r <= 12'hABA;
			12'h0E4 : dout_r <= 12'hABD;
			12'h0E5 : dout_r <= 12'hAC0;
			12'h0E6 : dout_r <= 12'hAC3;
			12'h0E7 : dout_r <= 12'hAC6;
			12'h0E8 : dout_r <= 12'hAC9;
			12'h0E9 : dout_r <= 12'hACC;
			12'h0EA : dout_r <= 12'hACF;
			12'h0EB : dout_r <= 12'hAD2;
			12'h0EC : dout_r <= 12'hAD4;
			12'h0ED : dout_r <= 12'hAD7;
			12'h0EE : dout_r <= 12'hADA;
			12'h0EF : dout_r <= 12'hADD;
			12'h0F0 : dout_r <= 12'hAE0;
			12'h0F1 : dout_r <= 12'hAE3;
			12'h0F2 : dout_r <= 12'hAE6;
			12'h0F3 : dout_r <= 12'hAE9;
			12'h0F4 : dout_r <= 12'hAEC;
			12'h0F5 : dout_r <= 12'hAEF;
			12'h0F6 : dout_r <= 12'hAF2;
			12'h0F7 : dout_r <= 12'hAF5;
			12'h0F8 : dout_r <= 12'hAF8;
			12'h0F9 : dout_r <= 12'hAFB;
			12'h0FA : dout_r <= 12'hAFD;
			12'h0FB : dout_r <= 12'hB00;
			12'h0FC : dout_r <= 12'hB03;
			12'h0FD : dout_r <= 12'hB06;
			12'h0FE : dout_r <= 12'hB09;
			12'h0FF : dout_r <= 12'hB0C;
			12'h100 : dout_r <= 12'hB0F;
			12'h101 : dout_r <= 12'hB12;
			12'h102 : dout_r <= 12'hB15;
			12'h103 : dout_r <= 12'hB18;
			12'h104 : dout_r <= 12'hB1A;
			12'h105 : dout_r <= 12'hB1D;
			12'h106 : dout_r <= 12'hB20;
			12'h107 : dout_r <= 12'hB23;
			12'h108 : dout_r <= 12'hB26;
			12'h109 : dout_r <= 12'hB29;
			12'h10A : dout_r <= 12'hB2C;
			12'h10B : dout_r <= 12'hB2F;
			12'h10C : dout_r <= 12'hB32;
			12'h10D : dout_r <= 12'hB34;
			12'h10E : dout_r <= 12'hB37;
			12'h10F : dout_r <= 12'hB3A;
			12'h110 : dout_r <= 12'hB3D;
			12'h111 : dout_r <= 12'hB40;
			12'h112 : dout_r <= 12'hB43;
			12'h113 : dout_r <= 12'hB46;
			12'h114 : dout_r <= 12'hB48;
			12'h115 : dout_r <= 12'hB4B;
			12'h116 : dout_r <= 12'hB4E;
			12'h117 : dout_r <= 12'hB51;
			12'h118 : dout_r <= 12'hB54;
			12'h119 : dout_r <= 12'hB57;
			12'h11A : dout_r <= 12'hB5A;
			12'h11B : dout_r <= 12'hB5C;
			12'h11C : dout_r <= 12'hB5F;
			12'h11D : dout_r <= 12'hB62;
			12'h11E : dout_r <= 12'hB65;
			12'h11F : dout_r <= 12'hB68;
			12'h120 : dout_r <= 12'hB6B;
			12'h121 : dout_r <= 12'hB6E;
			12'h122 : dout_r <= 12'hB70;
			12'h123 : dout_r <= 12'hB73;
			12'h124 : dout_r <= 12'hB76;
			12'h125 : dout_r <= 12'hB79;
			12'h126 : dout_r <= 12'hB7C;
			12'h127 : dout_r <= 12'hB7F;
			12'h128 : dout_r <= 12'hB81;
			12'h129 : dout_r <= 12'hB84;
			12'h12A : dout_r <= 12'hB87;
			12'h12B : dout_r <= 12'hB8A;
			12'h12C : dout_r <= 12'hB8D;
			12'h12D : dout_r <= 12'hB8F;
			12'h12E : dout_r <= 12'hB92;
			12'h12F : dout_r <= 12'hB95;
			12'h130 : dout_r <= 12'hB98;
			12'h131 : dout_r <= 12'hB9B;
			12'h132 : dout_r <= 12'hB9D;
			12'h133 : dout_r <= 12'hBA0;
			12'h134 : dout_r <= 12'hBA3;
			12'h135 : dout_r <= 12'hBA6;
			12'h136 : dout_r <= 12'hBA9;
			12'h137 : dout_r <= 12'hBAB;
			12'h138 : dout_r <= 12'hBAE;
			12'h139 : dout_r <= 12'hBB1;
			12'h13A : dout_r <= 12'hBB4;
			12'h13B : dout_r <= 12'hBB7;
			12'h13C : dout_r <= 12'hBB9;
			12'h13D : dout_r <= 12'hBBC;
			12'h13E : dout_r <= 12'hBBF;
			12'h13F : dout_r <= 12'hBC2;
			12'h140 : dout_r <= 12'hBC4;
			12'h141 : dout_r <= 12'hBC7;
			12'h142 : dout_r <= 12'hBCA;
			12'h143 : dout_r <= 12'hBCD;
			12'h144 : dout_r <= 12'hBD0;
			12'h145 : dout_r <= 12'hBD2;
			12'h146 : dout_r <= 12'hBD5;
			12'h147 : dout_r <= 12'hBD8;
			12'h148 : dout_r <= 12'hBDB;
			12'h149 : dout_r <= 12'hBDD;
			12'h14A : dout_r <= 12'hBE0;
			12'h14B : dout_r <= 12'hBE3;
			12'h14C : dout_r <= 12'hBE6;
			12'h14D : dout_r <= 12'hBE8;
			12'h14E : dout_r <= 12'hBEB;
			12'h14F : dout_r <= 12'hBEE;
			12'h150 : dout_r <= 12'hBF0;
			12'h151 : dout_r <= 12'hBF3;
			12'h152 : dout_r <= 12'hBF6;
			12'h153 : dout_r <= 12'hBF9;
			12'h154 : dout_r <= 12'hBFB;
			12'h155 : dout_r <= 12'hBFE;
			12'h156 : dout_r <= 12'hC01;
			12'h157 : dout_r <= 12'hC04;
			12'h158 : dout_r <= 12'hC06;
			12'h159 : dout_r <= 12'hC09;
			12'h15A : dout_r <= 12'hC0C;
			12'h15B : dout_r <= 12'hC0E;
			12'h15C : dout_r <= 12'hC11;
			12'h15D : dout_r <= 12'hC14;
			12'h15E : dout_r <= 12'hC16;
			12'h15F : dout_r <= 12'hC19;
			12'h160 : dout_r <= 12'hC1C;
			12'h161 : dout_r <= 12'hC1F;
			12'h162 : dout_r <= 12'hC21;
			12'h163 : dout_r <= 12'hC24;
			12'h164 : dout_r <= 12'hC27;
			12'h165 : dout_r <= 12'hC29;
			12'h166 : dout_r <= 12'hC2C;
			12'h167 : dout_r <= 12'hC2F;
			12'h168 : dout_r <= 12'hC31;
			12'h169 : dout_r <= 12'hC34;
			12'h16A : dout_r <= 12'hC37;
			12'h16B : dout_r <= 12'hC39;
			12'h16C : dout_r <= 12'hC3C;
			12'h16D : dout_r <= 12'hC3F;
			12'h16E : dout_r <= 12'hC41;
			12'h16F : dout_r <= 12'hC44;
			12'h170 : dout_r <= 12'hC47;
			12'h171 : dout_r <= 12'hC49;
			12'h172 : dout_r <= 12'hC4C;
			12'h173 : dout_r <= 12'hC4F;
			12'h174 : dout_r <= 12'hC51;
			12'h175 : dout_r <= 12'hC54;
			12'h176 : dout_r <= 12'hC57;
			12'h177 : dout_r <= 12'hC59;
			12'h178 : dout_r <= 12'hC5C;
			12'h179 : dout_r <= 12'hC5E;
			12'h17A : dout_r <= 12'hC61;
			12'h17B : dout_r <= 12'hC64;
			12'h17C : dout_r <= 12'hC66;
			12'h17D : dout_r <= 12'hC69;
			12'h17E : dout_r <= 12'hC6C;
			12'h17F : dout_r <= 12'hC6E;
			12'h180 : dout_r <= 12'hC71;
			12'h181 : dout_r <= 12'hC73;
			12'h182 : dout_r <= 12'hC76;
			12'h183 : dout_r <= 12'hC79;
			12'h184 : dout_r <= 12'hC7B;
			12'h185 : dout_r <= 12'hC7E;
			12'h186 : dout_r <= 12'hC80;
			12'h187 : dout_r <= 12'hC83;
			12'h188 : dout_r <= 12'hC86;
			12'h189 : dout_r <= 12'hC88;
			12'h18A : dout_r <= 12'hC8B;
			12'h18B : dout_r <= 12'hC8D;
			12'h18C : dout_r <= 12'hC90;
			12'h18D : dout_r <= 12'hC92;
			12'h18E : dout_r <= 12'hC95;
			12'h18F : dout_r <= 12'hC98;
			12'h190 : dout_r <= 12'hC9A;
			12'h191 : dout_r <= 12'hC9D;
			12'h192 : dout_r <= 12'hC9F;
			12'h193 : dout_r <= 12'hCA2;
			12'h194 : dout_r <= 12'hCA4;
			12'h195 : dout_r <= 12'hCA7;
			12'h196 : dout_r <= 12'hCAA;
			12'h197 : dout_r <= 12'hCAC;
			12'h198 : dout_r <= 12'hCAF;
			12'h199 : dout_r <= 12'hCB1;
			12'h19A : dout_r <= 12'hCB4;
			12'h19B : dout_r <= 12'hCB6;
			12'h19C : dout_r <= 12'hCB9;
			12'h19D : dout_r <= 12'hCBB;
			12'h19E : dout_r <= 12'hCBE;
			12'h19F : dout_r <= 12'hCC0;
			12'h1A0 : dout_r <= 12'hCC3;
			12'h1A1 : dout_r <= 12'hCC5;
			12'h1A2 : dout_r <= 12'hCC8;
			12'h1A3 : dout_r <= 12'hCCA;
			12'h1A4 : dout_r <= 12'hCCD;
			12'h1A5 : dout_r <= 12'hCCF;
			12'h1A6 : dout_r <= 12'hCD2;
			12'h1A7 : dout_r <= 12'hCD4;
			12'h1A8 : dout_r <= 12'hCD7;
			12'h1A9 : dout_r <= 12'hCD9;
			12'h1AA : dout_r <= 12'hCDC;
			12'h1AB : dout_r <= 12'hCDE;
			12'h1AC : dout_r <= 12'hCE1;
			12'h1AD : dout_r <= 12'hCE3;
			12'h1AE : dout_r <= 12'hCE6;
			12'h1AF : dout_r <= 12'hCE8;
			12'h1B0 : dout_r <= 12'hCEB;
			12'h1B1 : dout_r <= 12'hCED;
			12'h1B2 : dout_r <= 12'hCF0;
			12'h1B3 : dout_r <= 12'hCF2;
			12'h1B4 : dout_r <= 12'hCF5;
			12'h1B5 : dout_r <= 12'hCF7;
			12'h1B6 : dout_r <= 12'hCFA;
			12'h1B7 : dout_r <= 12'hCFC;
			12'h1B8 : dout_r <= 12'hCFF;
			12'h1B9 : dout_r <= 12'hD01;
			12'h1BA : dout_r <= 12'hD03;
			12'h1BB : dout_r <= 12'hD06;
			12'h1BC : dout_r <= 12'hD08;
			12'h1BD : dout_r <= 12'hD0B;
			12'h1BE : dout_r <= 12'hD0D;
			12'h1BF : dout_r <= 12'hD10;
			12'h1C0 : dout_r <= 12'hD12;
			12'h1C1 : dout_r <= 12'hD15;
			12'h1C2 : dout_r <= 12'hD17;
			12'h1C3 : dout_r <= 12'hD19;
			12'h1C4 : dout_r <= 12'hD1C;
			12'h1C5 : dout_r <= 12'hD1E;
			12'h1C6 : dout_r <= 12'hD21;
			12'h1C7 : dout_r <= 12'hD23;
			12'h1C8 : dout_r <= 12'hD25;
			12'h1C9 : dout_r <= 12'hD28;
			12'h1CA : dout_r <= 12'hD2A;
			12'h1CB : dout_r <= 12'hD2D;
			12'h1CC : dout_r <= 12'hD2F;
			12'h1CD : dout_r <= 12'hD31;
			12'h1CE : dout_r <= 12'hD34;
			12'h1CF : dout_r <= 12'hD36;
			12'h1D0 : dout_r <= 12'hD39;
			12'h1D1 : dout_r <= 12'hD3B;
			12'h1D2 : dout_r <= 12'hD3D;
			12'h1D3 : dout_r <= 12'hD40;
			12'h1D4 : dout_r <= 12'hD42;
			12'h1D5 : dout_r <= 12'hD44;
			12'h1D6 : dout_r <= 12'hD47;
			12'h1D7 : dout_r <= 12'hD49;
			12'h1D8 : dout_r <= 12'hD4B;
			12'h1D9 : dout_r <= 12'hD4E;
			12'h1DA : dout_r <= 12'hD50;
			12'h1DB : dout_r <= 12'hD53;
			12'h1DC : dout_r <= 12'hD55;
			12'h1DD : dout_r <= 12'hD57;
			12'h1DE : dout_r <= 12'hD5A;
			12'h1DF : dout_r <= 12'hD5C;
			12'h1E0 : dout_r <= 12'hD5E;
			12'h1E1 : dout_r <= 12'hD61;
			12'h1E2 : dout_r <= 12'hD63;
			12'h1E3 : dout_r <= 12'hD65;
			12'h1E4 : dout_r <= 12'hD67;
			12'h1E5 : dout_r <= 12'hD6A;
			12'h1E6 : dout_r <= 12'hD6C;
			12'h1E7 : dout_r <= 12'hD6E;
			12'h1E8 : dout_r <= 12'hD71;
			12'h1E9 : dout_r <= 12'hD73;
			12'h1EA : dout_r <= 12'hD75;
			12'h1EB : dout_r <= 12'hD78;
			12'h1EC : dout_r <= 12'hD7A;
			12'h1ED : dout_r <= 12'hD7C;
			12'h1EE : dout_r <= 12'hD7E;
			12'h1EF : dout_r <= 12'hD81;
			12'h1F0 : dout_r <= 12'hD83;
			12'h1F1 : dout_r <= 12'hD85;
			12'h1F2 : dout_r <= 12'hD88;
			12'h1F3 : dout_r <= 12'hD8A;
			12'h1F4 : dout_r <= 12'hD8C;
			12'h1F5 : dout_r <= 12'hD8E;
			12'h1F6 : dout_r <= 12'hD91;
			12'h1F7 : dout_r <= 12'hD93;
			12'h1F8 : dout_r <= 12'hD95;
			12'h1F9 : dout_r <= 12'hD97;
			12'h1FA : dout_r <= 12'hD9A;
			12'h1FB : dout_r <= 12'hD9C;
			12'h1FC : dout_r <= 12'hD9E;
			12'h1FD : dout_r <= 12'hDA0;
			12'h1FE : dout_r <= 12'hDA3;
			12'h1FF : dout_r <= 12'hDA5;
			12'h200 : dout_r <= 12'hDA7;
			12'h201 : dout_r <= 12'hDA9;
			12'h202 : dout_r <= 12'hDAB;
			12'h203 : dout_r <= 12'hDAE;
			12'h204 : dout_r <= 12'hDB0;
			12'h205 : dout_r <= 12'hDB2;
			12'h206 : dout_r <= 12'hDB4;
			12'h207 : dout_r <= 12'hDB6;
			12'h208 : dout_r <= 12'hDB9;
			12'h209 : dout_r <= 12'hDBB;
			12'h20A : dout_r <= 12'hDBD;
			12'h20B : dout_r <= 12'hDBF;
			12'h20C : dout_r <= 12'hDC1;
			12'h20D : dout_r <= 12'hDC4;
			12'h20E : dout_r <= 12'hDC6;
			12'h20F : dout_r <= 12'hDC8;
			12'h210 : dout_r <= 12'hDCA;
			12'h211 : dout_r <= 12'hDCC;
			12'h212 : dout_r <= 12'hDCE;
			12'h213 : dout_r <= 12'hDD1;
			12'h214 : dout_r <= 12'hDD3;
			12'h215 : dout_r <= 12'hDD5;
			12'h216 : dout_r <= 12'hDD7;
			12'h217 : dout_r <= 12'hDD9;
			12'h218 : dout_r <= 12'hDDB;
			12'h219 : dout_r <= 12'hDDD;
			12'h21A : dout_r <= 12'hDE0;
			12'h21B : dout_r <= 12'hDE2;
			12'h21C : dout_r <= 12'hDE4;
			12'h21D : dout_r <= 12'hDE6;
			12'h21E : dout_r <= 12'hDE8;
			12'h21F : dout_r <= 12'hDEA;
			12'h220 : dout_r <= 12'hDEC;
			12'h221 : dout_r <= 12'hDEE;
			12'h222 : dout_r <= 12'hDF0;
			12'h223 : dout_r <= 12'hDF3;
			12'h224 : dout_r <= 12'hDF5;
			12'h225 : dout_r <= 12'hDF7;
			12'h226 : dout_r <= 12'hDF9;
			12'h227 : dout_r <= 12'hDFB;
			12'h228 : dout_r <= 12'hDFD;
			12'h229 : dout_r <= 12'hDFF;
			12'h22A : dout_r <= 12'hE01;
			12'h22B : dout_r <= 12'hE03;
			12'h22C : dout_r <= 12'hE05;
			12'h22D : dout_r <= 12'hE07;
			12'h22E : dout_r <= 12'hE09;
			12'h22F : dout_r <= 12'hE0B;
			12'h230 : dout_r <= 12'hE0E;
			12'h231 : dout_r <= 12'hE10;
			12'h232 : dout_r <= 12'hE12;
			12'h233 : dout_r <= 12'hE14;
			12'h234 : dout_r <= 12'hE16;
			12'h235 : dout_r <= 12'hE18;
			12'h236 : dout_r <= 12'hE1A;
			12'h237 : dout_r <= 12'hE1C;
			12'h238 : dout_r <= 12'hE1E;
			12'h239 : dout_r <= 12'hE20;
			12'h23A : dout_r <= 12'hE22;
			12'h23B : dout_r <= 12'hE24;
			12'h23C : dout_r <= 12'hE26;
			12'h23D : dout_r <= 12'hE28;
			12'h23E : dout_r <= 12'hE2A;
			12'h23F : dout_r <= 12'hE2C;
			12'h240 : dout_r <= 12'hE2E;
			12'h241 : dout_r <= 12'hE30;
			12'h242 : dout_r <= 12'hE32;
			12'h243 : dout_r <= 12'hE34;
			12'h244 : dout_r <= 12'hE36;
			12'h245 : dout_r <= 12'hE38;
			12'h246 : dout_r <= 12'hE3A;
			12'h247 : dout_r <= 12'hE3C;
			12'h248 : dout_r <= 12'hE3E;
			12'h249 : dout_r <= 12'hE40;
			12'h24A : dout_r <= 12'hE42;
			12'h24B : dout_r <= 12'hE44;
			12'h24C : dout_r <= 12'hE45;
			12'h24D : dout_r <= 12'hE47;
			12'h24E : dout_r <= 12'hE49;
			12'h24F : dout_r <= 12'hE4B;
			12'h250 : dout_r <= 12'hE4D;
			12'h251 : dout_r <= 12'hE4F;
			12'h252 : dout_r <= 12'hE51;
			12'h253 : dout_r <= 12'hE53;
			12'h254 : dout_r <= 12'hE55;
			12'h255 : dout_r <= 12'hE57;
			12'h256 : dout_r <= 12'hE59;
			12'h257 : dout_r <= 12'hE5B;
			12'h258 : dout_r <= 12'hE5D;
			12'h259 : dout_r <= 12'hE5E;
			12'h25A : dout_r <= 12'hE60;
			12'h25B : dout_r <= 12'hE62;
			12'h25C : dout_r <= 12'hE64;
			12'h25D : dout_r <= 12'hE66;
			12'h25E : dout_r <= 12'hE68;
			12'h25F : dout_r <= 12'hE6A;
			12'h260 : dout_r <= 12'hE6C;
			12'h261 : dout_r <= 12'hE6E;
			12'h262 : dout_r <= 12'hE6F;
			12'h263 : dout_r <= 12'hE71;
			12'h264 : dout_r <= 12'hE73;
			12'h265 : dout_r <= 12'hE75;
			12'h266 : dout_r <= 12'hE77;
			12'h267 : dout_r <= 12'hE79;
			12'h268 : dout_r <= 12'hE7B;
			12'h269 : dout_r <= 12'hE7C;
			12'h26A : dout_r <= 12'hE7E;
			12'h26B : dout_r <= 12'hE80;
			12'h26C : dout_r <= 12'hE82;
			12'h26D : dout_r <= 12'hE84;
			12'h26E : dout_r <= 12'hE85;
			12'h26F : dout_r <= 12'hE87;
			12'h270 : dout_r <= 12'hE89;
			12'h271 : dout_r <= 12'hE8B;
			12'h272 : dout_r <= 12'hE8D;
			12'h273 : dout_r <= 12'hE8F;
			12'h274 : dout_r <= 12'hE90;
			12'h275 : dout_r <= 12'hE92;
			12'h276 : dout_r <= 12'hE94;
			12'h277 : dout_r <= 12'hE96;
			12'h278 : dout_r <= 12'hE97;
			12'h279 : dout_r <= 12'hE99;
			12'h27A : dout_r <= 12'hE9B;
			12'h27B : dout_r <= 12'hE9D;
			12'h27C : dout_r <= 12'hE9F;
			12'h27D : dout_r <= 12'hEA0;
			12'h27E : dout_r <= 12'hEA2;
			12'h27F : dout_r <= 12'hEA4;
			12'h280 : dout_r <= 12'hEA6;
			12'h281 : dout_r <= 12'hEA7;
			12'h282 : dout_r <= 12'hEA9;
			12'h283 : dout_r <= 12'hEAB;
			12'h284 : dout_r <= 12'hEAC;
			12'h285 : dout_r <= 12'hEAE;
			12'h286 : dout_r <= 12'hEB0;
			12'h287 : dout_r <= 12'hEB2;
			12'h288 : dout_r <= 12'hEB3;
			12'h289 : dout_r <= 12'hEB5;
			12'h28A : dout_r <= 12'hEB7;
			12'h28B : dout_r <= 12'hEB8;
			12'h28C : dout_r <= 12'hEBA;
			12'h28D : dout_r <= 12'hEBC;
			12'h28E : dout_r <= 12'hEBE;
			12'h28F : dout_r <= 12'hEBF;
			12'h290 : dout_r <= 12'hEC1;
			12'h291 : dout_r <= 12'hEC3;
			12'h292 : dout_r <= 12'hEC4;
			12'h293 : dout_r <= 12'hEC6;
			12'h294 : dout_r <= 12'hEC8;
			12'h295 : dout_r <= 12'hEC9;
			12'h296 : dout_r <= 12'hECB;
			12'h297 : dout_r <= 12'hECD;
			12'h298 : dout_r <= 12'hECE;
			12'h299 : dout_r <= 12'hED0;
			12'h29A : dout_r <= 12'hED2;
			12'h29B : dout_r <= 12'hED3;
			12'h29C : dout_r <= 12'hED5;
			12'h29D : dout_r <= 12'hED6;
			12'h29E : dout_r <= 12'hED8;
			12'h29F : dout_r <= 12'hEDA;
			12'h2A0 : dout_r <= 12'hEDB;
			12'h2A1 : dout_r <= 12'hEDD;
			12'h2A2 : dout_r <= 12'hEDE;
			12'h2A3 : dout_r <= 12'hEE0;
			12'h2A4 : dout_r <= 12'hEE2;
			12'h2A5 : dout_r <= 12'hEE3;
			12'h2A6 : dout_r <= 12'hEE5;
			12'h2A7 : dout_r <= 12'hEE6;
			12'h2A8 : dout_r <= 12'hEE8;
			12'h2A9 : dout_r <= 12'hEEA;
			12'h2AA : dout_r <= 12'hEEB;
			12'h2AB : dout_r <= 12'hEED;
			12'h2AC : dout_r <= 12'hEEE;
			12'h2AD : dout_r <= 12'hEF0;
			12'h2AE : dout_r <= 12'hEF1;
			12'h2AF : dout_r <= 12'hEF3;
			12'h2B0 : dout_r <= 12'hEF5;
			12'h2B1 : dout_r <= 12'hEF6;
			12'h2B2 : dout_r <= 12'hEF8;
			12'h2B3 : dout_r <= 12'hEF9;
			12'h2B4 : dout_r <= 12'hEFB;
			12'h2B5 : dout_r <= 12'hEFC;
			12'h2B6 : dout_r <= 12'hEFE;
			12'h2B7 : dout_r <= 12'hEFF;
			12'h2B8 : dout_r <= 12'hF01;
			12'h2B9 : dout_r <= 12'hF02;
			12'h2BA : dout_r <= 12'hF04;
			12'h2BB : dout_r <= 12'hF05;
			12'h2BC : dout_r <= 12'hF07;
			12'h2BD : dout_r <= 12'hF08;
			12'h2BE : dout_r <= 12'hF0A;
			12'h2BF : dout_r <= 12'hF0B;
			12'h2C0 : dout_r <= 12'hF0D;
			12'h2C1 : dout_r <= 12'hF0E;
			12'h2C2 : dout_r <= 12'hF10;
			12'h2C3 : dout_r <= 12'hF11;
			12'h2C4 : dout_r <= 12'hF13;
			12'h2C5 : dout_r <= 12'hF14;
			12'h2C6 : dout_r <= 12'hF16;
			12'h2C7 : dout_r <= 12'hF17;
			12'h2C8 : dout_r <= 12'hF18;
			12'h2C9 : dout_r <= 12'hF1A;
			12'h2CA : dout_r <= 12'hF1B;
			12'h2CB : dout_r <= 12'hF1D;
			12'h2CC : dout_r <= 12'hF1E;
			12'h2CD : dout_r <= 12'hF20;
			12'h2CE : dout_r <= 12'hF21;
			12'h2CF : dout_r <= 12'hF23;
			12'h2D0 : dout_r <= 12'hF24;
			12'h2D1 : dout_r <= 12'hF25;
			12'h2D2 : dout_r <= 12'hF27;
			12'h2D3 : dout_r <= 12'hF28;
			12'h2D4 : dout_r <= 12'hF2A;
			12'h2D5 : dout_r <= 12'hF2B;
			12'h2D6 : dout_r <= 12'hF2C;
			12'h2D7 : dout_r <= 12'hF2E;
			12'h2D8 : dout_r <= 12'hF2F;
			12'h2D9 : dout_r <= 12'hF30;
			12'h2DA : dout_r <= 12'hF32;
			12'h2DB : dout_r <= 12'hF33;
			12'h2DC : dout_r <= 12'hF35;
			12'h2DD : dout_r <= 12'hF36;
			12'h2DE : dout_r <= 12'hF37;
			12'h2DF : dout_r <= 12'hF39;
			12'h2E0 : dout_r <= 12'hF3A;
			12'h2E1 : dout_r <= 12'hF3B;
			12'h2E2 : dout_r <= 12'hF3D;
			12'h2E3 : dout_r <= 12'hF3E;
			12'h2E4 : dout_r <= 12'hF3F;
			12'h2E5 : dout_r <= 12'hF41;
			12'h2E6 : dout_r <= 12'hF42;
			12'h2E7 : dout_r <= 12'hF43;
			12'h2E8 : dout_r <= 12'hF45;
			12'h2E9 : dout_r <= 12'hF46;
			12'h2EA : dout_r <= 12'hF47;
			12'h2EB : dout_r <= 12'hF48;
			12'h2EC : dout_r <= 12'hF4A;
			12'h2ED : dout_r <= 12'hF4B;
			12'h2EE : dout_r <= 12'hF4C;
			12'h2EF : dout_r <= 12'hF4E;
			12'h2F0 : dout_r <= 12'hF4F;
			12'h2F1 : dout_r <= 12'hF50;
			12'h2F2 : dout_r <= 12'hF51;
			12'h2F3 : dout_r <= 12'hF53;
			12'h2F4 : dout_r <= 12'hF54;
			12'h2F5 : dout_r <= 12'hF55;
			12'h2F6 : dout_r <= 12'hF56;
			12'h2F7 : dout_r <= 12'hF58;
			12'h2F8 : dout_r <= 12'hF59;
			12'h2F9 : dout_r <= 12'hF5A;
			12'h2FA : dout_r <= 12'hF5B;
			12'h2FB : dout_r <= 12'hF5D;
			12'h2FC : dout_r <= 12'hF5E;
			12'h2FD : dout_r <= 12'hF5F;
			12'h2FE : dout_r <= 12'hF60;
			12'h2FF : dout_r <= 12'hF61;
			12'h300 : dout_r <= 12'hF63;
			12'h301 : dout_r <= 12'hF64;
			12'h302 : dout_r <= 12'hF65;
			12'h303 : dout_r <= 12'hF66;
			12'h304 : dout_r <= 12'hF67;
			12'h305 : dout_r <= 12'hF69;
			12'h306 : dout_r <= 12'hF6A;
			12'h307 : dout_r <= 12'hF6B;
			12'h308 : dout_r <= 12'hF6C;
			12'h309 : dout_r <= 12'hF6D;
			12'h30A : dout_r <= 12'hF6E;
			12'h30B : dout_r <= 12'hF70;
			12'h30C : dout_r <= 12'hF71;
			12'h30D : dout_r <= 12'hF72;
			12'h30E : dout_r <= 12'hF73;
			12'h30F : dout_r <= 12'hF74;
			12'h310 : dout_r <= 12'hF75;
			12'h311 : dout_r <= 12'hF76;
			12'h312 : dout_r <= 12'hF78;
			12'h313 : dout_r <= 12'hF79;
			12'h314 : dout_r <= 12'hF7A;
			12'h315 : dout_r <= 12'hF7B;
			12'h316 : dout_r <= 12'hF7C;
			12'h317 : dout_r <= 12'hF7D;
			12'h318 : dout_r <= 12'hF7E;
			12'h319 : dout_r <= 12'hF7F;
			12'h31A : dout_r <= 12'hF80;
			12'h31B : dout_r <= 12'hF81;
			12'h31C : dout_r <= 12'hF83;
			12'h31D : dout_r <= 12'hF84;
			12'h31E : dout_r <= 12'hF85;
			12'h31F : dout_r <= 12'hF86;
			12'h320 : dout_r <= 12'hF87;
			12'h321 : dout_r <= 12'hF88;
			12'h322 : dout_r <= 12'hF89;
			12'h323 : dout_r <= 12'hF8A;
			12'h324 : dout_r <= 12'hF8B;
			12'h325 : dout_r <= 12'hF8C;
			12'h326 : dout_r <= 12'hF8D;
			12'h327 : dout_r <= 12'hF8E;
			12'h328 : dout_r <= 12'hF8F;
			12'h329 : dout_r <= 12'hF90;
			12'h32A : dout_r <= 12'hF91;
			12'h32B : dout_r <= 12'hF92;
			12'h32C : dout_r <= 12'hF93;
			12'h32D : dout_r <= 12'hF94;
			12'h32E : dout_r <= 12'hF95;
			12'h32F : dout_r <= 12'hF96;
			12'h330 : dout_r <= 12'hF97;
			12'h331 : dout_r <= 12'hF98;
			12'h332 : dout_r <= 12'hF99;
			12'h333 : dout_r <= 12'hF9A;
			12'h334 : dout_r <= 12'hF9B;
			12'h335 : dout_r <= 12'hF9C;
			12'h336 : dout_r <= 12'hF9D;
			12'h337 : dout_r <= 12'hF9E;
			12'h338 : dout_r <= 12'hF9F;
			12'h339 : dout_r <= 12'hFA0;
			12'h33A : dout_r <= 12'hFA1;
			12'h33B : dout_r <= 12'hFA2;
			12'h33C : dout_r <= 12'hFA3;
			12'h33D : dout_r <= 12'hFA4;
			12'h33E : dout_r <= 12'hFA5;
			12'h33F : dout_r <= 12'hFA5;
			12'h340 : dout_r <= 12'hFA6;
			12'h341 : dout_r <= 12'hFA7;
			12'h342 : dout_r <= 12'hFA8;
			12'h343 : dout_r <= 12'hFA9;
			12'h344 : dout_r <= 12'hFAA;
			12'h345 : dout_r <= 12'hFAB;
			12'h346 : dout_r <= 12'hFAC;
			12'h347 : dout_r <= 12'hFAD;
			12'h348 : dout_r <= 12'hFAE;
			12'h349 : dout_r <= 12'hFAE;
			12'h34A : dout_r <= 12'hFAF;
			12'h34B : dout_r <= 12'hFB0;
			12'h34C : dout_r <= 12'hFB1;
			12'h34D : dout_r <= 12'hFB2;
			12'h34E : dout_r <= 12'hFB3;
			12'h34F : dout_r <= 12'hFB4;
			12'h350 : dout_r <= 12'hFB4;
			12'h351 : dout_r <= 12'hFB5;
			12'h352 : dout_r <= 12'hFB6;
			12'h353 : dout_r <= 12'hFB7;
			12'h354 : dout_r <= 12'hFB8;
			12'h355 : dout_r <= 12'hFB8;
			12'h356 : dout_r <= 12'hFB9;
			12'h357 : dout_r <= 12'hFBA;
			12'h358 : dout_r <= 12'hFBB;
			12'h359 : dout_r <= 12'hFBC;
			12'h35A : dout_r <= 12'hFBC;
			12'h35B : dout_r <= 12'hFBD;
			12'h35C : dout_r <= 12'hFBE;
			12'h35D : dout_r <= 12'hFBF;
			12'h35E : dout_r <= 12'hFC0;
			12'h35F : dout_r <= 12'hFC0;
			12'h360 : dout_r <= 12'hFC1;
			12'h361 : dout_r <= 12'hFC2;
			12'h362 : dout_r <= 12'hFC3;
			12'h363 : dout_r <= 12'hFC3;
			12'h364 : dout_r <= 12'hFC4;
			12'h365 : dout_r <= 12'hFC5;
			12'h366 : dout_r <= 12'hFC6;
			12'h367 : dout_r <= 12'hFC6;
			12'h368 : dout_r <= 12'hFC7;
			12'h369 : dout_r <= 12'hFC8;
			12'h36A : dout_r <= 12'hFC9;
			12'h36B : dout_r <= 12'hFC9;
			12'h36C : dout_r <= 12'hFCA;
			12'h36D : dout_r <= 12'hFCB;
			12'h36E : dout_r <= 12'hFCB;
			12'h36F : dout_r <= 12'hFCC;
			12'h370 : dout_r <= 12'hFCD;
			12'h371 : dout_r <= 12'hFCD;
			12'h372 : dout_r <= 12'hFCE;
			12'h373 : dout_r <= 12'hFCF;
			12'h374 : dout_r <= 12'hFCF;
			12'h375 : dout_r <= 12'hFD0;
			12'h376 : dout_r <= 12'hFD1;
			12'h377 : dout_r <= 12'hFD1;
			12'h378 : dout_r <= 12'hFD2;
			12'h379 : dout_r <= 12'hFD3;
			12'h37A : dout_r <= 12'hFD3;
			12'h37B : dout_r <= 12'hFD4;
			12'h37C : dout_r <= 12'hFD5;
			12'h37D : dout_r <= 12'hFD5;
			12'h37E : dout_r <= 12'hFD6;
			12'h37F : dout_r <= 12'hFD7;
			12'h380 : dout_r <= 12'hFD7;
			12'h381 : dout_r <= 12'hFD8;
			12'h382 : dout_r <= 12'hFD8;
			12'h383 : dout_r <= 12'hFD9;
			12'h384 : dout_r <= 12'hFDA;
			12'h385 : dout_r <= 12'hFDA;
			12'h386 : dout_r <= 12'hFDB;
			12'h387 : dout_r <= 12'hFDB;
			12'h388 : dout_r <= 12'hFDC;
			12'h389 : dout_r <= 12'hFDC;
			12'h38A : dout_r <= 12'hFDD;
			12'h38B : dout_r <= 12'hFDE;
			12'h38C : dout_r <= 12'hFDE;
			12'h38D : dout_r <= 12'hFDF;
			12'h38E : dout_r <= 12'hFDF;
			12'h38F : dout_r <= 12'hFE0;
			12'h390 : dout_r <= 12'hFE0;
			12'h391 : dout_r <= 12'hFE1;
			12'h392 : dout_r <= 12'hFE1;
			12'h393 : dout_r <= 12'hFE2;
			12'h394 : dout_r <= 12'hFE2;
			12'h395 : dout_r <= 12'hFE3;
			12'h396 : dout_r <= 12'hFE3;
			12'h397 : dout_r <= 12'hFE4;
			12'h398 : dout_r <= 12'hFE5;
			12'h399 : dout_r <= 12'hFE5;
			12'h39A : dout_r <= 12'hFE5;
			12'h39B : dout_r <= 12'hFE6;
			12'h39C : dout_r <= 12'hFE6;
			12'h39D : dout_r <= 12'hFE7;
			12'h39E : dout_r <= 12'hFE7;
			12'h39F : dout_r <= 12'hFE8;
			12'h3A0 : dout_r <= 12'hFE8;
			12'h3A1 : dout_r <= 12'hFE9;
			12'h3A2 : dout_r <= 12'hFE9;
			12'h3A3 : dout_r <= 12'hFEA;
			12'h3A4 : dout_r <= 12'hFEA;
			12'h3A5 : dout_r <= 12'hFEB;
			12'h3A6 : dout_r <= 12'hFEB;
			12'h3A7 : dout_r <= 12'hFEB;
			12'h3A8 : dout_r <= 12'hFEC;
			12'h3A9 : dout_r <= 12'hFEC;
			12'h3AA : dout_r <= 12'hFED;
			12'h3AB : dout_r <= 12'hFED;
			12'h3AC : dout_r <= 12'hFEE;
			12'h3AD : dout_r <= 12'hFEE;
			12'h3AE : dout_r <= 12'hFEE;
			12'h3AF : dout_r <= 12'hFEF;
			12'h3B0 : dout_r <= 12'hFEF;
			12'h3B1 : dout_r <= 12'hFEF;
			12'h3B2 : dout_r <= 12'hFF0;
			12'h3B3 : dout_r <= 12'hFF0;
			12'h3B4 : dout_r <= 12'hFF1;
			12'h3B5 : dout_r <= 12'hFF1;
			12'h3B6 : dout_r <= 12'hFF1;
			12'h3B7 : dout_r <= 12'hFF2;
			12'h3B8 : dout_r <= 12'hFF2;
			12'h3B9 : dout_r <= 12'hFF2;
			12'h3BA : dout_r <= 12'hFF3;
			12'h3BB : dout_r <= 12'hFF3;
			12'h3BC : dout_r <= 12'hFF3;
			12'h3BD : dout_r <= 12'hFF4;
			12'h3BE : dout_r <= 12'hFF4;
			12'h3BF : dout_r <= 12'hFF4;
			12'h3C0 : dout_r <= 12'hFF5;
			12'h3C1 : dout_r <= 12'hFF5;
			12'h3C2 : dout_r <= 12'hFF5;
			12'h3C3 : dout_r <= 12'hFF6;
			12'h3C4 : dout_r <= 12'hFF6;
			12'h3C5 : dout_r <= 12'hFF6;
			12'h3C6 : dout_r <= 12'hFF6;
			12'h3C7 : dout_r <= 12'hFF7;
			12'h3C8 : dout_r <= 12'hFF7;
			12'h3C9 : dout_r <= 12'hFF7;
			12'h3CA : dout_r <= 12'hFF7;
			12'h3CB : dout_r <= 12'hFF8;
			12'h3CC : dout_r <= 12'hFF8;
			12'h3CD : dout_r <= 12'hFF8;
			12'h3CE : dout_r <= 12'hFF8;
			12'h3CF : dout_r <= 12'hFF9;
			12'h3D0 : dout_r <= 12'hFF9;
			12'h3D1 : dout_r <= 12'hFF9;
			12'h3D2 : dout_r <= 12'hFF9;
			12'h3D3 : dout_r <= 12'hFFA;
			12'h3D4 : dout_r <= 12'hFFA;
			12'h3D5 : dout_r <= 12'hFFA;
			12'h3D6 : dout_r <= 12'hFFA;
			12'h3D7 : dout_r <= 12'hFFA;
			12'h3D8 : dout_r <= 12'hFFB;
			12'h3D9 : dout_r <= 12'hFFB;
			12'h3DA : dout_r <= 12'hFFB;
			12'h3DB : dout_r <= 12'hFFB;
			12'h3DC : dout_r <= 12'hFFB;
			12'h3DD : dout_r <= 12'hFFC;
			12'h3DE : dout_r <= 12'hFFC;
			12'h3DF : dout_r <= 12'hFFC;
			12'h3E0 : dout_r <= 12'hFFC;
			12'h3E1 : dout_r <= 12'hFFC;
			12'h3E2 : dout_r <= 12'hFFC;
			12'h3E3 : dout_r <= 12'hFFC;
			12'h3E4 : dout_r <= 12'hFFD;
			12'h3E5 : dout_r <= 12'hFFD;
			12'h3E6 : dout_r <= 12'hFFD;
			12'h3E7 : dout_r <= 12'hFFD;
			12'h3E8 : dout_r <= 12'hFFD;
			12'h3E9 : dout_r <= 12'hFFD;
			12'h3EA : dout_r <= 12'hFFD;
			12'h3EB : dout_r <= 12'hFFD;
			12'h3EC : dout_r <= 12'hFFE;
			12'h3ED : dout_r <= 12'hFFE;
			12'h3EE : dout_r <= 12'hFFE;
			12'h3EF : dout_r <= 12'hFFE;
			12'h3F0 : dout_r <= 12'hFFE;
			12'h3F1 : dout_r <= 12'hFFE;
			12'h3F2 : dout_r <= 12'hFFE;
			12'h3F3 : dout_r <= 12'hFFE;
			12'h3F4 : dout_r <= 12'hFFE;
			12'h3F5 : dout_r <= 12'hFFE;
			12'h3F6 : dout_r <= 12'hFFE;
			12'h3F7 : dout_r <= 12'hFFE;
			12'h3F8 : dout_r <= 12'hFFE;
			12'h3F9 : dout_r <= 12'hFFE;
			12'h3FA : dout_r <= 12'hFFE;
			12'h3FB : dout_r <= 12'hFFE;
			12'h3FC : dout_r <= 12'hFFE;
			12'h3FD : dout_r <= 12'hFFE;
			12'h3FE : dout_r <= 12'hFFE;
			12'h3FF : dout_r <= 12'hFFE;
			12'h400 : dout_r <= 12'hFFF;
			12'h401 : dout_r <= 12'hFFE;
			12'h402 : dout_r <= 12'hFFE;
			12'h403 : dout_r <= 12'hFFE;
			12'h404 : dout_r <= 12'hFFE;
			12'h405 : dout_r <= 12'hFFE;
			12'h406 : dout_r <= 12'hFFE;
			12'h407 : dout_r <= 12'hFFE;
			12'h408 : dout_r <= 12'hFFE;
			12'h409 : dout_r <= 12'hFFE;
			12'h40A : dout_r <= 12'hFFE;
			12'h40B : dout_r <= 12'hFFE;
			12'h40C : dout_r <= 12'hFFE;
			12'h40D : dout_r <= 12'hFFE;
			12'h40E : dout_r <= 12'hFFE;
			12'h40F : dout_r <= 12'hFFE;
			12'h410 : dout_r <= 12'hFFE;
			12'h411 : dout_r <= 12'hFFE;
			12'h412 : dout_r <= 12'hFFE;
			12'h413 : dout_r <= 12'hFFE;
			12'h414 : dout_r <= 12'hFFE;
			12'h415 : dout_r <= 12'hFFD;
			12'h416 : dout_r <= 12'hFFD;
			12'h417 : dout_r <= 12'hFFD;
			12'h418 : dout_r <= 12'hFFD;
			12'h419 : dout_r <= 12'hFFD;
			12'h41A : dout_r <= 12'hFFD;
			12'h41B : dout_r <= 12'hFFD;
			12'h41C : dout_r <= 12'hFFD;
			12'h41D : dout_r <= 12'hFFC;
			12'h41E : dout_r <= 12'hFFC;
			12'h41F : dout_r <= 12'hFFC;
			12'h420 : dout_r <= 12'hFFC;
			12'h421 : dout_r <= 12'hFFC;
			12'h422 : dout_r <= 12'hFFC;
			12'h423 : dout_r <= 12'hFFC;
			12'h424 : dout_r <= 12'hFFB;
			12'h425 : dout_r <= 12'hFFB;
			12'h426 : dout_r <= 12'hFFB;
			12'h427 : dout_r <= 12'hFFB;
			12'h428 : dout_r <= 12'hFFB;
			12'h429 : dout_r <= 12'hFFA;
			12'h42A : dout_r <= 12'hFFA;
			12'h42B : dout_r <= 12'hFFA;
			12'h42C : dout_r <= 12'hFFA;
			12'h42D : dout_r <= 12'hFFA;
			12'h42E : dout_r <= 12'hFF9;
			12'h42F : dout_r <= 12'hFF9;
			12'h430 : dout_r <= 12'hFF9;
			12'h431 : dout_r <= 12'hFF9;
			12'h432 : dout_r <= 12'hFF8;
			12'h433 : dout_r <= 12'hFF8;
			12'h434 : dout_r <= 12'hFF8;
			12'h435 : dout_r <= 12'hFF8;
			12'h436 : dout_r <= 12'hFF7;
			12'h437 : dout_r <= 12'hFF7;
			12'h438 : dout_r <= 12'hFF7;
			12'h439 : dout_r <= 12'hFF7;
			12'h43A : dout_r <= 12'hFF6;
			12'h43B : dout_r <= 12'hFF6;
			12'h43C : dout_r <= 12'hFF6;
			12'h43D : dout_r <= 12'hFF6;
			12'h43E : dout_r <= 12'hFF5;
			12'h43F : dout_r <= 12'hFF5;
			12'h440 : dout_r <= 12'hFF5;
			12'h441 : dout_r <= 12'hFF4;
			12'h442 : dout_r <= 12'hFF4;
			12'h443 : dout_r <= 12'hFF4;
			12'h444 : dout_r <= 12'hFF3;
			12'h445 : dout_r <= 12'hFF3;
			12'h446 : dout_r <= 12'hFF3;
			12'h447 : dout_r <= 12'hFF2;
			12'h448 : dout_r <= 12'hFF2;
			12'h449 : dout_r <= 12'hFF2;
			12'h44A : dout_r <= 12'hFF1;
			12'h44B : dout_r <= 12'hFF1;
			12'h44C : dout_r <= 12'hFF1;
			12'h44D : dout_r <= 12'hFF0;
			12'h44E : dout_r <= 12'hFF0;
			12'h44F : dout_r <= 12'hFEF;
			12'h450 : dout_r <= 12'hFEF;
			12'h451 : dout_r <= 12'hFEF;
			12'h452 : dout_r <= 12'hFEE;
			12'h453 : dout_r <= 12'hFEE;
			12'h454 : dout_r <= 12'hFEE;
			12'h455 : dout_r <= 12'hFED;
			12'h456 : dout_r <= 12'hFED;
			12'h457 : dout_r <= 12'hFEC;
			12'h458 : dout_r <= 12'hFEC;
			12'h459 : dout_r <= 12'hFEB;
			12'h45A : dout_r <= 12'hFEB;
			12'h45B : dout_r <= 12'hFEB;
			12'h45C : dout_r <= 12'hFEA;
			12'h45D : dout_r <= 12'hFEA;
			12'h45E : dout_r <= 12'hFE9;
			12'h45F : dout_r <= 12'hFE9;
			12'h460 : dout_r <= 12'hFE8;
			12'h461 : dout_r <= 12'hFE8;
			12'h462 : dout_r <= 12'hFE7;
			12'h463 : dout_r <= 12'hFE7;
			12'h464 : dout_r <= 12'hFE6;
			12'h465 : dout_r <= 12'hFE6;
			12'h466 : dout_r <= 12'hFE5;
			12'h467 : dout_r <= 12'hFE5;
			12'h468 : dout_r <= 12'hFE5;
			12'h469 : dout_r <= 12'hFE4;
			12'h46A : dout_r <= 12'hFE3;
			12'h46B : dout_r <= 12'hFE3;
			12'h46C : dout_r <= 12'hFE2;
			12'h46D : dout_r <= 12'hFE2;
			12'h46E : dout_r <= 12'hFE1;
			12'h46F : dout_r <= 12'hFE1;
			12'h470 : dout_r <= 12'hFE0;
			12'h471 : dout_r <= 12'hFE0;
			12'h472 : dout_r <= 12'hFDF;
			12'h473 : dout_r <= 12'hFDF;
			12'h474 : dout_r <= 12'hFDE;
			12'h475 : dout_r <= 12'hFDE;
			12'h476 : dout_r <= 12'hFDD;
			12'h477 : dout_r <= 12'hFDC;
			12'h478 : dout_r <= 12'hFDC;
			12'h479 : dout_r <= 12'hFDB;
			12'h47A : dout_r <= 12'hFDB;
			12'h47B : dout_r <= 12'hFDA;
			12'h47C : dout_r <= 12'hFDA;
			12'h47D : dout_r <= 12'hFD9;
			12'h47E : dout_r <= 12'hFD8;
			12'h47F : dout_r <= 12'hFD8;
			12'h480 : dout_r <= 12'hFD7;
			12'h481 : dout_r <= 12'hFD7;
			12'h482 : dout_r <= 12'hFD6;
			12'h483 : dout_r <= 12'hFD5;
			12'h484 : dout_r <= 12'hFD5;
			12'h485 : dout_r <= 12'hFD4;
			12'h486 : dout_r <= 12'hFD3;
			12'h487 : dout_r <= 12'hFD3;
			12'h488 : dout_r <= 12'hFD2;
			12'h489 : dout_r <= 12'hFD1;
			12'h48A : dout_r <= 12'hFD1;
			12'h48B : dout_r <= 12'hFD0;
			12'h48C : dout_r <= 12'hFCF;
			12'h48D : dout_r <= 12'hFCF;
			12'h48E : dout_r <= 12'hFCE;
			12'h48F : dout_r <= 12'hFCD;
			12'h490 : dout_r <= 12'hFCD;
			12'h491 : dout_r <= 12'hFCC;
			12'h492 : dout_r <= 12'hFCB;
			12'h493 : dout_r <= 12'hFCB;
			12'h494 : dout_r <= 12'hFCA;
			12'h495 : dout_r <= 12'hFC9;
			12'h496 : dout_r <= 12'hFC9;
			12'h497 : dout_r <= 12'hFC8;
			12'h498 : dout_r <= 12'hFC7;
			12'h499 : dout_r <= 12'hFC6;
			12'h49A : dout_r <= 12'hFC6;
			12'h49B : dout_r <= 12'hFC5;
			12'h49C : dout_r <= 12'hFC4;
			12'h49D : dout_r <= 12'hFC3;
			12'h49E : dout_r <= 12'hFC3;
			12'h49F : dout_r <= 12'hFC2;
			12'h4A0 : dout_r <= 12'hFC1;
			12'h4A1 : dout_r <= 12'hFC0;
			12'h4A2 : dout_r <= 12'hFC0;
			12'h4A3 : dout_r <= 12'hFBF;
			12'h4A4 : dout_r <= 12'hFBE;
			12'h4A5 : dout_r <= 12'hFBD;
			12'h4A6 : dout_r <= 12'hFBC;
			12'h4A7 : dout_r <= 12'hFBC;
			12'h4A8 : dout_r <= 12'hFBB;
			12'h4A9 : dout_r <= 12'hFBA;
			12'h4AA : dout_r <= 12'hFB9;
			12'h4AB : dout_r <= 12'hFB8;
			12'h4AC : dout_r <= 12'hFB8;
			12'h4AD : dout_r <= 12'hFB7;
			12'h4AE : dout_r <= 12'hFB6;
			12'h4AF : dout_r <= 12'hFB5;
			12'h4B0 : dout_r <= 12'hFB4;
			12'h4B1 : dout_r <= 12'hFB4;
			12'h4B2 : dout_r <= 12'hFB3;
			12'h4B3 : dout_r <= 12'hFB2;
			12'h4B4 : dout_r <= 12'hFB1;
			12'h4B5 : dout_r <= 12'hFB0;
			12'h4B6 : dout_r <= 12'hFAF;
			12'h4B7 : dout_r <= 12'hFAE;
			12'h4B8 : dout_r <= 12'hFAE;
			12'h4B9 : dout_r <= 12'hFAD;
			12'h4BA : dout_r <= 12'hFAC;
			12'h4BB : dout_r <= 12'hFAB;
			12'h4BC : dout_r <= 12'hFAA;
			12'h4BD : dout_r <= 12'hFA9;
			12'h4BE : dout_r <= 12'hFA8;
			12'h4BF : dout_r <= 12'hFA7;
			12'h4C0 : dout_r <= 12'hFA6;
			12'h4C1 : dout_r <= 12'hFA5;
			12'h4C2 : dout_r <= 12'hFA5;
			12'h4C3 : dout_r <= 12'hFA4;
			12'h4C4 : dout_r <= 12'hFA3;
			12'h4C5 : dout_r <= 12'hFA2;
			12'h4C6 : dout_r <= 12'hFA1;
			12'h4C7 : dout_r <= 12'hFA0;
			12'h4C8 : dout_r <= 12'hF9F;
			12'h4C9 : dout_r <= 12'hF9E;
			12'h4CA : dout_r <= 12'hF9D;
			12'h4CB : dout_r <= 12'hF9C;
			12'h4CC : dout_r <= 12'hF9B;
			12'h4CD : dout_r <= 12'hF9A;
			12'h4CE : dout_r <= 12'hF99;
			12'h4CF : dout_r <= 12'hF98;
			12'h4D0 : dout_r <= 12'hF97;
			12'h4D1 : dout_r <= 12'hF96;
			12'h4D2 : dout_r <= 12'hF95;
			12'h4D3 : dout_r <= 12'hF94;
			12'h4D4 : dout_r <= 12'hF93;
			12'h4D5 : dout_r <= 12'hF92;
			12'h4D6 : dout_r <= 12'hF91;
			12'h4D7 : dout_r <= 12'hF90;
			12'h4D8 : dout_r <= 12'hF8F;
			12'h4D9 : dout_r <= 12'hF8E;
			12'h4DA : dout_r <= 12'hF8D;
			12'h4DB : dout_r <= 12'hF8C;
			12'h4DC : dout_r <= 12'hF8B;
			12'h4DD : dout_r <= 12'hF8A;
			12'h4DE : dout_r <= 12'hF89;
			12'h4DF : dout_r <= 12'hF88;
			12'h4E0 : dout_r <= 12'hF87;
			12'h4E1 : dout_r <= 12'hF86;
			12'h4E2 : dout_r <= 12'hF85;
			12'h4E3 : dout_r <= 12'hF84;
			12'h4E4 : dout_r <= 12'hF83;
			12'h4E5 : dout_r <= 12'hF81;
			12'h4E6 : dout_r <= 12'hF80;
			12'h4E7 : dout_r <= 12'hF7F;
			12'h4E8 : dout_r <= 12'hF7E;
			12'h4E9 : dout_r <= 12'hF7D;
			12'h4EA : dout_r <= 12'hF7C;
			12'h4EB : dout_r <= 12'hF7B;
			12'h4EC : dout_r <= 12'hF7A;
			12'h4ED : dout_r <= 12'hF79;
			12'h4EE : dout_r <= 12'hF78;
			12'h4EF : dout_r <= 12'hF76;
			12'h4F0 : dout_r <= 12'hF75;
			12'h4F1 : dout_r <= 12'hF74;
			12'h4F2 : dout_r <= 12'hF73;
			12'h4F3 : dout_r <= 12'hF72;
			12'h4F4 : dout_r <= 12'hF71;
			12'h4F5 : dout_r <= 12'hF70;
			12'h4F6 : dout_r <= 12'hF6E;
			12'h4F7 : dout_r <= 12'hF6D;
			12'h4F8 : dout_r <= 12'hF6C;
			12'h4F9 : dout_r <= 12'hF6B;
			12'h4FA : dout_r <= 12'hF6A;
			12'h4FB : dout_r <= 12'hF69;
			12'h4FC : dout_r <= 12'hF67;
			12'h4FD : dout_r <= 12'hF66;
			12'h4FE : dout_r <= 12'hF65;
			12'h4FF : dout_r <= 12'hF64;
			12'h500 : dout_r <= 12'hF63;
			12'h501 : dout_r <= 12'hF61;
			12'h502 : dout_r <= 12'hF60;
			12'h503 : dout_r <= 12'hF5F;
			12'h504 : dout_r <= 12'hF5E;
			12'h505 : dout_r <= 12'hF5D;
			12'h506 : dout_r <= 12'hF5B;
			12'h507 : dout_r <= 12'hF5A;
			12'h508 : dout_r <= 12'hF59;
			12'h509 : dout_r <= 12'hF58;
			12'h50A : dout_r <= 12'hF56;
			12'h50B : dout_r <= 12'hF55;
			12'h50C : dout_r <= 12'hF54;
			12'h50D : dout_r <= 12'hF53;
			12'h50E : dout_r <= 12'hF51;
			12'h50F : dout_r <= 12'hF50;
			12'h510 : dout_r <= 12'hF4F;
			12'h511 : dout_r <= 12'hF4E;
			12'h512 : dout_r <= 12'hF4C;
			12'h513 : dout_r <= 12'hF4B;
			12'h514 : dout_r <= 12'hF4A;
			12'h515 : dout_r <= 12'hF48;
			12'h516 : dout_r <= 12'hF47;
			12'h517 : dout_r <= 12'hF46;
			12'h518 : dout_r <= 12'hF45;
			12'h519 : dout_r <= 12'hF43;
			12'h51A : dout_r <= 12'hF42;
			12'h51B : dout_r <= 12'hF41;
			12'h51C : dout_r <= 12'hF3F;
			12'h51D : dout_r <= 12'hF3E;
			12'h51E : dout_r <= 12'hF3D;
			12'h51F : dout_r <= 12'hF3B;
			12'h520 : dout_r <= 12'hF3A;
			12'h521 : dout_r <= 12'hF39;
			12'h522 : dout_r <= 12'hF37;
			12'h523 : dout_r <= 12'hF36;
			12'h524 : dout_r <= 12'hF35;
			12'h525 : dout_r <= 12'hF33;
			12'h526 : dout_r <= 12'hF32;
			12'h527 : dout_r <= 12'hF30;
			12'h528 : dout_r <= 12'hF2F;
			12'h529 : dout_r <= 12'hF2E;
			12'h52A : dout_r <= 12'hF2C;
			12'h52B : dout_r <= 12'hF2B;
			12'h52C : dout_r <= 12'hF2A;
			12'h52D : dout_r <= 12'hF28;
			12'h52E : dout_r <= 12'hF27;
			12'h52F : dout_r <= 12'hF25;
			12'h530 : dout_r <= 12'hF24;
			12'h531 : dout_r <= 12'hF23;
			12'h532 : dout_r <= 12'hF21;
			12'h533 : dout_r <= 12'hF20;
			12'h534 : dout_r <= 12'hF1E;
			12'h535 : dout_r <= 12'hF1D;
			12'h536 : dout_r <= 12'hF1B;
			12'h537 : dout_r <= 12'hF1A;
			12'h538 : dout_r <= 12'hF18;
			12'h539 : dout_r <= 12'hF17;
			12'h53A : dout_r <= 12'hF16;
			12'h53B : dout_r <= 12'hF14;
			12'h53C : dout_r <= 12'hF13;
			12'h53D : dout_r <= 12'hF11;
			12'h53E : dout_r <= 12'hF10;
			12'h53F : dout_r <= 12'hF0E;
			12'h540 : dout_r <= 12'hF0D;
			12'h541 : dout_r <= 12'hF0B;
			12'h542 : dout_r <= 12'hF0A;
			12'h543 : dout_r <= 12'hF08;
			12'h544 : dout_r <= 12'hF07;
			12'h545 : dout_r <= 12'hF05;
			12'h546 : dout_r <= 12'hF04;
			12'h547 : dout_r <= 12'hF02;
			12'h548 : dout_r <= 12'hF01;
			12'h549 : dout_r <= 12'hEFF;
			12'h54A : dout_r <= 12'hEFE;
			12'h54B : dout_r <= 12'hEFC;
			12'h54C : dout_r <= 12'hEFB;
			12'h54D : dout_r <= 12'hEF9;
			12'h54E : dout_r <= 12'hEF8;
			12'h54F : dout_r <= 12'hEF6;
			12'h550 : dout_r <= 12'hEF5;
			12'h551 : dout_r <= 12'hEF3;
			12'h552 : dout_r <= 12'hEF1;
			12'h553 : dout_r <= 12'hEF0;
			12'h554 : dout_r <= 12'hEEE;
			12'h555 : dout_r <= 12'hEED;
			12'h556 : dout_r <= 12'hEEB;
			12'h557 : dout_r <= 12'hEEA;
			12'h558 : dout_r <= 12'hEE8;
			12'h559 : dout_r <= 12'hEE6;
			12'h55A : dout_r <= 12'hEE5;
			12'h55B : dout_r <= 12'hEE3;
			12'h55C : dout_r <= 12'hEE2;
			12'h55D : dout_r <= 12'hEE0;
			12'h55E : dout_r <= 12'hEDE;
			12'h55F : dout_r <= 12'hEDD;
			12'h560 : dout_r <= 12'hEDB;
			12'h561 : dout_r <= 12'hEDA;
			12'h562 : dout_r <= 12'hED8;
			12'h563 : dout_r <= 12'hED6;
			12'h564 : dout_r <= 12'hED5;
			12'h565 : dout_r <= 12'hED3;
			12'h566 : dout_r <= 12'hED2;
			12'h567 : dout_r <= 12'hED0;
			12'h568 : dout_r <= 12'hECE;
			12'h569 : dout_r <= 12'hECD;
			12'h56A : dout_r <= 12'hECB;
			12'h56B : dout_r <= 12'hEC9;
			12'h56C : dout_r <= 12'hEC8;
			12'h56D : dout_r <= 12'hEC6;
			12'h56E : dout_r <= 12'hEC4;
			12'h56F : dout_r <= 12'hEC3;
			12'h570 : dout_r <= 12'hEC1;
			12'h571 : dout_r <= 12'hEBF;
			12'h572 : dout_r <= 12'hEBE;
			12'h573 : dout_r <= 12'hEBC;
			12'h574 : dout_r <= 12'hEBA;
			12'h575 : dout_r <= 12'hEB8;
			12'h576 : dout_r <= 12'hEB7;
			12'h577 : dout_r <= 12'hEB5;
			12'h578 : dout_r <= 12'hEB3;
			12'h579 : dout_r <= 12'hEB2;
			12'h57A : dout_r <= 12'hEB0;
			12'h57B : dout_r <= 12'hEAE;
			12'h57C : dout_r <= 12'hEAC;
			12'h57D : dout_r <= 12'hEAB;
			12'h57E : dout_r <= 12'hEA9;
			12'h57F : dout_r <= 12'hEA7;
			12'h580 : dout_r <= 12'hEA6;
			12'h581 : dout_r <= 12'hEA4;
			12'h582 : dout_r <= 12'hEA2;
			12'h583 : dout_r <= 12'hEA0;
			12'h584 : dout_r <= 12'hE9F;
			12'h585 : dout_r <= 12'hE9D;
			12'h586 : dout_r <= 12'hE9B;
			12'h587 : dout_r <= 12'hE99;
			12'h588 : dout_r <= 12'hE97;
			12'h589 : dout_r <= 12'hE96;
			12'h58A : dout_r <= 12'hE94;
			12'h58B : dout_r <= 12'hE92;
			12'h58C : dout_r <= 12'hE90;
			12'h58D : dout_r <= 12'hE8F;
			12'h58E : dout_r <= 12'hE8D;
			12'h58F : dout_r <= 12'hE8B;
			12'h590 : dout_r <= 12'hE89;
			12'h591 : dout_r <= 12'hE87;
			12'h592 : dout_r <= 12'hE85;
			12'h593 : dout_r <= 12'hE84;
			12'h594 : dout_r <= 12'hE82;
			12'h595 : dout_r <= 12'hE80;
			12'h596 : dout_r <= 12'hE7E;
			12'h597 : dout_r <= 12'hE7C;
			12'h598 : dout_r <= 12'hE7B;
			12'h599 : dout_r <= 12'hE79;
			12'h59A : dout_r <= 12'hE77;
			12'h59B : dout_r <= 12'hE75;
			12'h59C : dout_r <= 12'hE73;
			12'h59D : dout_r <= 12'hE71;
			12'h59E : dout_r <= 12'hE6F;
			12'h59F : dout_r <= 12'hE6E;
			12'h5A0 : dout_r <= 12'hE6C;
			12'h5A1 : dout_r <= 12'hE6A;
			12'h5A2 : dout_r <= 12'hE68;
			12'h5A3 : dout_r <= 12'hE66;
			12'h5A4 : dout_r <= 12'hE64;
			12'h5A5 : dout_r <= 12'hE62;
			12'h5A6 : dout_r <= 12'hE60;
			12'h5A7 : dout_r <= 12'hE5E;
			12'h5A8 : dout_r <= 12'hE5D;
			12'h5A9 : dout_r <= 12'hE5B;
			12'h5AA : dout_r <= 12'hE59;
			12'h5AB : dout_r <= 12'hE57;
			12'h5AC : dout_r <= 12'hE55;
			12'h5AD : dout_r <= 12'hE53;
			12'h5AE : dout_r <= 12'hE51;
			12'h5AF : dout_r <= 12'hE4F;
			12'h5B0 : dout_r <= 12'hE4D;
			12'h5B1 : dout_r <= 12'hE4B;
			12'h5B2 : dout_r <= 12'hE49;
			12'h5B3 : dout_r <= 12'hE47;
			12'h5B4 : dout_r <= 12'hE45;
			12'h5B5 : dout_r <= 12'hE44;
			12'h5B6 : dout_r <= 12'hE42;
			12'h5B7 : dout_r <= 12'hE40;
			12'h5B8 : dout_r <= 12'hE3E;
			12'h5B9 : dout_r <= 12'hE3C;
			12'h5BA : dout_r <= 12'hE3A;
			12'h5BB : dout_r <= 12'hE38;
			12'h5BC : dout_r <= 12'hE36;
			12'h5BD : dout_r <= 12'hE34;
			12'h5BE : dout_r <= 12'hE32;
			12'h5BF : dout_r <= 12'hE30;
			12'h5C0 : dout_r <= 12'hE2E;
			12'h5C1 : dout_r <= 12'hE2C;
			12'h5C2 : dout_r <= 12'hE2A;
			12'h5C3 : dout_r <= 12'hE28;
			12'h5C4 : dout_r <= 12'hE26;
			12'h5C5 : dout_r <= 12'hE24;
			12'h5C6 : dout_r <= 12'hE22;
			12'h5C7 : dout_r <= 12'hE20;
			12'h5C8 : dout_r <= 12'hE1E;
			12'h5C9 : dout_r <= 12'hE1C;
			12'h5CA : dout_r <= 12'hE1A;
			12'h5CB : dout_r <= 12'hE18;
			12'h5CC : dout_r <= 12'hE16;
			12'h5CD : dout_r <= 12'hE14;
			12'h5CE : dout_r <= 12'hE12;
			12'h5CF : dout_r <= 12'hE10;
			12'h5D0 : dout_r <= 12'hE0E;
			12'h5D1 : dout_r <= 12'hE0B;
			12'h5D2 : dout_r <= 12'hE09;
			12'h5D3 : dout_r <= 12'hE07;
			12'h5D4 : dout_r <= 12'hE05;
			12'h5D5 : dout_r <= 12'hE03;
			12'h5D6 : dout_r <= 12'hE01;
			12'h5D7 : dout_r <= 12'hDFF;
			12'h5D8 : dout_r <= 12'hDFD;
			12'h5D9 : dout_r <= 12'hDFB;
			12'h5DA : dout_r <= 12'hDF9;
			12'h5DB : dout_r <= 12'hDF7;
			12'h5DC : dout_r <= 12'hDF5;
			12'h5DD : dout_r <= 12'hDF3;
			12'h5DE : dout_r <= 12'hDF0;
			12'h5DF : dout_r <= 12'hDEE;
			12'h5E0 : dout_r <= 12'hDEC;
			12'h5E1 : dout_r <= 12'hDEA;
			12'h5E2 : dout_r <= 12'hDE8;
			12'h5E3 : dout_r <= 12'hDE6;
			12'h5E4 : dout_r <= 12'hDE4;
			12'h5E5 : dout_r <= 12'hDE2;
			12'h5E6 : dout_r <= 12'hDE0;
			12'h5E7 : dout_r <= 12'hDDD;
			12'h5E8 : dout_r <= 12'hDDB;
			12'h5E9 : dout_r <= 12'hDD9;
			12'h5EA : dout_r <= 12'hDD7;
			12'h5EB : dout_r <= 12'hDD5;
			12'h5EC : dout_r <= 12'hDD3;
			12'h5ED : dout_r <= 12'hDD1;
			12'h5EE : dout_r <= 12'hDCE;
			12'h5EF : dout_r <= 12'hDCC;
			12'h5F0 : dout_r <= 12'hDCA;
			12'h5F1 : dout_r <= 12'hDC8;
			12'h5F2 : dout_r <= 12'hDC6;
			12'h5F3 : dout_r <= 12'hDC4;
			12'h5F4 : dout_r <= 12'hDC1;
			12'h5F5 : dout_r <= 12'hDBF;
			12'h5F6 : dout_r <= 12'hDBD;
			12'h5F7 : dout_r <= 12'hDBB;
			12'h5F8 : dout_r <= 12'hDB9;
			12'h5F9 : dout_r <= 12'hDB6;
			12'h5FA : dout_r <= 12'hDB4;
			12'h5FB : dout_r <= 12'hDB2;
			12'h5FC : dout_r <= 12'hDB0;
			12'h5FD : dout_r <= 12'hDAE;
			12'h5FE : dout_r <= 12'hDAB;
			12'h5FF : dout_r <= 12'hDA9;
			12'h600 : dout_r <= 12'hDA7;
			12'h601 : dout_r <= 12'hDA5;
			12'h602 : dout_r <= 12'hDA3;
			12'h603 : dout_r <= 12'hDA0;
			12'h604 : dout_r <= 12'hD9E;
			12'h605 : dout_r <= 12'hD9C;
			12'h606 : dout_r <= 12'hD9A;
			12'h607 : dout_r <= 12'hD97;
			12'h608 : dout_r <= 12'hD95;
			12'h609 : dout_r <= 12'hD93;
			12'h60A : dout_r <= 12'hD91;
			12'h60B : dout_r <= 12'hD8E;
			12'h60C : dout_r <= 12'hD8C;
			12'h60D : dout_r <= 12'hD8A;
			12'h60E : dout_r <= 12'hD88;
			12'h60F : dout_r <= 12'hD85;
			12'h610 : dout_r <= 12'hD83;
			12'h611 : dout_r <= 12'hD81;
			12'h612 : dout_r <= 12'hD7E;
			12'h613 : dout_r <= 12'hD7C;
			12'h614 : dout_r <= 12'hD7A;
			12'h615 : dout_r <= 12'hD78;
			12'h616 : dout_r <= 12'hD75;
			12'h617 : dout_r <= 12'hD73;
			12'h618 : dout_r <= 12'hD71;
			12'h619 : dout_r <= 12'hD6E;
			12'h61A : dout_r <= 12'hD6C;
			12'h61B : dout_r <= 12'hD6A;
			12'h61C : dout_r <= 12'hD67;
			12'h61D : dout_r <= 12'hD65;
			12'h61E : dout_r <= 12'hD63;
			12'h61F : dout_r <= 12'hD61;
			12'h620 : dout_r <= 12'hD5E;
			12'h621 : dout_r <= 12'hD5C;
			12'h622 : dout_r <= 12'hD5A;
			12'h623 : dout_r <= 12'hD57;
			12'h624 : dout_r <= 12'hD55;
			12'h625 : dout_r <= 12'hD53;
			12'h626 : dout_r <= 12'hD50;
			12'h627 : dout_r <= 12'hD4E;
			12'h628 : dout_r <= 12'hD4B;
			12'h629 : dout_r <= 12'hD49;
			12'h62A : dout_r <= 12'hD47;
			12'h62B : dout_r <= 12'hD44;
			12'h62C : dout_r <= 12'hD42;
			12'h62D : dout_r <= 12'hD40;
			12'h62E : dout_r <= 12'hD3D;
			12'h62F : dout_r <= 12'hD3B;
			12'h630 : dout_r <= 12'hD39;
			12'h631 : dout_r <= 12'hD36;
			12'h632 : dout_r <= 12'hD34;
			12'h633 : dout_r <= 12'hD31;
			12'h634 : dout_r <= 12'hD2F;
			12'h635 : dout_r <= 12'hD2D;
			12'h636 : dout_r <= 12'hD2A;
			12'h637 : dout_r <= 12'hD28;
			12'h638 : dout_r <= 12'hD25;
			12'h639 : dout_r <= 12'hD23;
			12'h63A : dout_r <= 12'hD21;
			12'h63B : dout_r <= 12'hD1E;
			12'h63C : dout_r <= 12'hD1C;
			12'h63D : dout_r <= 12'hD19;
			12'h63E : dout_r <= 12'hD17;
			12'h63F : dout_r <= 12'hD15;
			12'h640 : dout_r <= 12'hD12;
			12'h641 : dout_r <= 12'hD10;
			12'h642 : dout_r <= 12'hD0D;
			12'h643 : dout_r <= 12'hD0B;
			12'h644 : dout_r <= 12'hD08;
			12'h645 : dout_r <= 12'hD06;
			12'h646 : dout_r <= 12'hD03;
			12'h647 : dout_r <= 12'hD01;
			12'h648 : dout_r <= 12'hCFF;
			12'h649 : dout_r <= 12'hCFC;
			12'h64A : dout_r <= 12'hCFA;
			12'h64B : dout_r <= 12'hCF7;
			12'h64C : dout_r <= 12'hCF5;
			12'h64D : dout_r <= 12'hCF2;
			12'h64E : dout_r <= 12'hCF0;
			12'h64F : dout_r <= 12'hCED;
			12'h650 : dout_r <= 12'hCEB;
			12'h651 : dout_r <= 12'hCE8;
			12'h652 : dout_r <= 12'hCE6;
			12'h653 : dout_r <= 12'hCE3;
			12'h654 : dout_r <= 12'hCE1;
			12'h655 : dout_r <= 12'hCDE;
			12'h656 : dout_r <= 12'hCDC;
			12'h657 : dout_r <= 12'hCD9;
			12'h658 : dout_r <= 12'hCD7;
			12'h659 : dout_r <= 12'hCD4;
			12'h65A : dout_r <= 12'hCD2;
			12'h65B : dout_r <= 12'hCCF;
			12'h65C : dout_r <= 12'hCCD;
			12'h65D : dout_r <= 12'hCCA;
			12'h65E : dout_r <= 12'hCC8;
			12'h65F : dout_r <= 12'hCC5;
			12'h660 : dout_r <= 12'hCC3;
			12'h661 : dout_r <= 12'hCC0;
			12'h662 : dout_r <= 12'hCBE;
			12'h663 : dout_r <= 12'hCBB;
			12'h664 : dout_r <= 12'hCB9;
			12'h665 : dout_r <= 12'hCB6;
			12'h666 : dout_r <= 12'hCB4;
			12'h667 : dout_r <= 12'hCB1;
			12'h668 : dout_r <= 12'hCAF;
			12'h669 : dout_r <= 12'hCAC;
			12'h66A : dout_r <= 12'hCAA;
			12'h66B : dout_r <= 12'hCA7;
			12'h66C : dout_r <= 12'hCA4;
			12'h66D : dout_r <= 12'hCA2;
			12'h66E : dout_r <= 12'hC9F;
			12'h66F : dout_r <= 12'hC9D;
			12'h670 : dout_r <= 12'hC9A;
			12'h671 : dout_r <= 12'hC98;
			12'h672 : dout_r <= 12'hC95;
			12'h673 : dout_r <= 12'hC92;
			12'h674 : dout_r <= 12'hC90;
			12'h675 : dout_r <= 12'hC8D;
			12'h676 : dout_r <= 12'hC8B;
			12'h677 : dout_r <= 12'hC88;
			12'h678 : dout_r <= 12'hC86;
			12'h679 : dout_r <= 12'hC83;
			12'h67A : dout_r <= 12'hC80;
			12'h67B : dout_r <= 12'hC7E;
			12'h67C : dout_r <= 12'hC7B;
			12'h67D : dout_r <= 12'hC79;
			12'h67E : dout_r <= 12'hC76;
			12'h67F : dout_r <= 12'hC73;
			12'h680 : dout_r <= 12'hC71;
			12'h681 : dout_r <= 12'hC6E;
			12'h682 : dout_r <= 12'hC6C;
			12'h683 : dout_r <= 12'hC69;
			12'h684 : dout_r <= 12'hC66;
			12'h685 : dout_r <= 12'hC64;
			12'h686 : dout_r <= 12'hC61;
			12'h687 : dout_r <= 12'hC5E;
			12'h688 : dout_r <= 12'hC5C;
			12'h689 : dout_r <= 12'hC59;
			12'h68A : dout_r <= 12'hC57;
			12'h68B : dout_r <= 12'hC54;
			12'h68C : dout_r <= 12'hC51;
			12'h68D : dout_r <= 12'hC4F;
			12'h68E : dout_r <= 12'hC4C;
			12'h68F : dout_r <= 12'hC49;
			12'h690 : dout_r <= 12'hC47;
			12'h691 : dout_r <= 12'hC44;
			12'h692 : dout_r <= 12'hC41;
			12'h693 : dout_r <= 12'hC3F;
			12'h694 : dout_r <= 12'hC3C;
			12'h695 : dout_r <= 12'hC39;
			12'h696 : dout_r <= 12'hC37;
			12'h697 : dout_r <= 12'hC34;
			12'h698 : dout_r <= 12'hC31;
			12'h699 : dout_r <= 12'hC2F;
			12'h69A : dout_r <= 12'hC2C;
			12'h69B : dout_r <= 12'hC29;
			12'h69C : dout_r <= 12'hC27;
			12'h69D : dout_r <= 12'hC24;
			12'h69E : dout_r <= 12'hC21;
			12'h69F : dout_r <= 12'hC1F;
			12'h6A0 : dout_r <= 12'hC1C;
			12'h6A1 : dout_r <= 12'hC19;
			12'h6A2 : dout_r <= 12'hC16;
			12'h6A3 : dout_r <= 12'hC14;
			12'h6A4 : dout_r <= 12'hC11;
			12'h6A5 : dout_r <= 12'hC0E;
			12'h6A6 : dout_r <= 12'hC0C;
			12'h6A7 : dout_r <= 12'hC09;
			12'h6A8 : dout_r <= 12'hC06;
			12'h6A9 : dout_r <= 12'hC04;
			12'h6AA : dout_r <= 12'hC01;
			12'h6AB : dout_r <= 12'hBFE;
			12'h6AC : dout_r <= 12'hBFB;
			12'h6AD : dout_r <= 12'hBF9;
			12'h6AE : dout_r <= 12'hBF6;
			12'h6AF : dout_r <= 12'hBF3;
			12'h6B0 : dout_r <= 12'hBF0;
			12'h6B1 : dout_r <= 12'hBEE;
			12'h6B2 : dout_r <= 12'hBEB;
			12'h6B3 : dout_r <= 12'hBE8;
			12'h6B4 : dout_r <= 12'hBE6;
			12'h6B5 : dout_r <= 12'hBE3;
			12'h6B6 : dout_r <= 12'hBE0;
			12'h6B7 : dout_r <= 12'hBDD;
			12'h6B8 : dout_r <= 12'hBDB;
			12'h6B9 : dout_r <= 12'hBD8;
			12'h6BA : dout_r <= 12'hBD5;
			12'h6BB : dout_r <= 12'hBD2;
			12'h6BC : dout_r <= 12'hBD0;
			12'h6BD : dout_r <= 12'hBCD;
			12'h6BE : dout_r <= 12'hBCA;
			12'h6BF : dout_r <= 12'hBC7;
			12'h6C0 : dout_r <= 12'hBC4;
			12'h6C1 : dout_r <= 12'hBC2;
			12'h6C2 : dout_r <= 12'hBBF;
			12'h6C3 : dout_r <= 12'hBBC;
			12'h6C4 : dout_r <= 12'hBB9;
			12'h6C5 : dout_r <= 12'hBB7;
			12'h6C6 : dout_r <= 12'hBB4;
			12'h6C7 : dout_r <= 12'hBB1;
			12'h6C8 : dout_r <= 12'hBAE;
			12'h6C9 : dout_r <= 12'hBAB;
			12'h6CA : dout_r <= 12'hBA9;
			12'h6CB : dout_r <= 12'hBA6;
			12'h6CC : dout_r <= 12'hBA3;
			12'h6CD : dout_r <= 12'hBA0;
			12'h6CE : dout_r <= 12'hB9D;
			12'h6CF : dout_r <= 12'hB9B;
			12'h6D0 : dout_r <= 12'hB98;
			12'h6D1 : dout_r <= 12'hB95;
			12'h6D2 : dout_r <= 12'hB92;
			12'h6D3 : dout_r <= 12'hB8F;
			12'h6D4 : dout_r <= 12'hB8D;
			12'h6D5 : dout_r <= 12'hB8A;
			12'h6D6 : dout_r <= 12'hB87;
			12'h6D7 : dout_r <= 12'hB84;
			12'h6D8 : dout_r <= 12'hB81;
			12'h6D9 : dout_r <= 12'hB7F;
			12'h6DA : dout_r <= 12'hB7C;
			12'h6DB : dout_r <= 12'hB79;
			12'h6DC : dout_r <= 12'hB76;
			12'h6DD : dout_r <= 12'hB73;
			12'h6DE : dout_r <= 12'hB70;
			12'h6DF : dout_r <= 12'hB6E;
			12'h6E0 : dout_r <= 12'hB6B;
			12'h6E1 : dout_r <= 12'hB68;
			12'h6E2 : dout_r <= 12'hB65;
			12'h6E3 : dout_r <= 12'hB62;
			12'h6E4 : dout_r <= 12'hB5F;
			12'h6E5 : dout_r <= 12'hB5C;
			12'h6E6 : dout_r <= 12'hB5A;
			12'h6E7 : dout_r <= 12'hB57;
			12'h6E8 : dout_r <= 12'hB54;
			12'h6E9 : dout_r <= 12'hB51;
			12'h6EA : dout_r <= 12'hB4E;
			12'h6EB : dout_r <= 12'hB4B;
			12'h6EC : dout_r <= 12'hB48;
			12'h6ED : dout_r <= 12'hB46;
			12'h6EE : dout_r <= 12'hB43;
			12'h6EF : dout_r <= 12'hB40;
			12'h6F0 : dout_r <= 12'hB3D;
			12'h6F1 : dout_r <= 12'hB3A;
			12'h6F2 : dout_r <= 12'hB37;
			12'h6F3 : dout_r <= 12'hB34;
			12'h6F4 : dout_r <= 12'hB32;
			12'h6F5 : dout_r <= 12'hB2F;
			12'h6F6 : dout_r <= 12'hB2C;
			12'h6F7 : dout_r <= 12'hB29;
			12'h6F8 : dout_r <= 12'hB26;
			12'h6F9 : dout_r <= 12'hB23;
			12'h6FA : dout_r <= 12'hB20;
			12'h6FB : dout_r <= 12'hB1D;
			12'h6FC : dout_r <= 12'hB1A;
			12'h6FD : dout_r <= 12'hB18;
			12'h6FE : dout_r <= 12'hB15;
			12'h6FF : dout_r <= 12'hB12;
			12'h700 : dout_r <= 12'hB0F;
			12'h701 : dout_r <= 12'hB0C;
			12'h702 : dout_r <= 12'hB09;
			12'h703 : dout_r <= 12'hB06;
			12'h704 : dout_r <= 12'hB03;
			12'h705 : dout_r <= 12'hB00;
			12'h706 : dout_r <= 12'hAFD;
			12'h707 : dout_r <= 12'hAFB;
			12'h708 : dout_r <= 12'hAF8;
			12'h709 : dout_r <= 12'hAF5;
			12'h70A : dout_r <= 12'hAF2;
			12'h70B : dout_r <= 12'hAEF;
			12'h70C : dout_r <= 12'hAEC;
			12'h70D : dout_r <= 12'hAE9;
			12'h70E : dout_r <= 12'hAE6;
			12'h70F : dout_r <= 12'hAE3;
			12'h710 : dout_r <= 12'hAE0;
			12'h711 : dout_r <= 12'hADD;
			12'h712 : dout_r <= 12'hADA;
			12'h713 : dout_r <= 12'hAD7;
			12'h714 : dout_r <= 12'hAD4;
			12'h715 : dout_r <= 12'hAD2;
			12'h716 : dout_r <= 12'hACF;
			12'h717 : dout_r <= 12'hACC;
			12'h718 : dout_r <= 12'hAC9;
			12'h719 : dout_r <= 12'hAC6;
			12'h71A : dout_r <= 12'hAC3;
			12'h71B : dout_r <= 12'hAC0;
			12'h71C : dout_r <= 12'hABD;
			12'h71D : dout_r <= 12'hABA;
			12'h71E : dout_r <= 12'hAB7;
			12'h71F : dout_r <= 12'hAB4;
			12'h720 : dout_r <= 12'hAB1;
			12'h721 : dout_r <= 12'hAAE;
			12'h722 : dout_r <= 12'hAAB;
			12'h723 : dout_r <= 12'hAA8;
			12'h724 : dout_r <= 12'hAA5;
			12'h725 : dout_r <= 12'hAA2;
			12'h726 : dout_r <= 12'hA9F;
			12'h727 : dout_r <= 12'hA9C;
			12'h728 : dout_r <= 12'hA99;
			12'h729 : dout_r <= 12'hA96;
			12'h72A : dout_r <= 12'hA93;
			12'h72B : dout_r <= 12'hA90;
			12'h72C : dout_r <= 12'hA8E;
			12'h72D : dout_r <= 12'hA8B;
			12'h72E : dout_r <= 12'hA88;
			12'h72F : dout_r <= 12'hA85;
			12'h730 : dout_r <= 12'hA82;
			12'h731 : dout_r <= 12'hA7F;
			12'h732 : dout_r <= 12'hA7C;
			12'h733 : dout_r <= 12'hA79;
			12'h734 : dout_r <= 12'hA76;
			12'h735 : dout_r <= 12'hA73;
			12'h736 : dout_r <= 12'hA70;
			12'h737 : dout_r <= 12'hA6D;
			12'h738 : dout_r <= 12'hA6A;
			12'h739 : dout_r <= 12'hA67;
			12'h73A : dout_r <= 12'hA64;
			12'h73B : dout_r <= 12'hA61;
			12'h73C : dout_r <= 12'hA5E;
			12'h73D : dout_r <= 12'hA5B;
			12'h73E : dout_r <= 12'hA58;
			12'h73F : dout_r <= 12'hA55;
			12'h740 : dout_r <= 12'hA52;
			12'h741 : dout_r <= 12'hA4F;
			12'h742 : dout_r <= 12'hA4C;
			12'h743 : dout_r <= 12'hA49;
			12'h744 : dout_r <= 12'hA46;
			12'h745 : dout_r <= 12'hA43;
			12'h746 : dout_r <= 12'hA40;
			12'h747 : dout_r <= 12'hA3D;
			12'h748 : dout_r <= 12'hA3A;
			12'h749 : dout_r <= 12'hA37;
			12'h74A : dout_r <= 12'hA34;
			12'h74B : dout_r <= 12'hA31;
			12'h74C : dout_r <= 12'hA2E;
			12'h74D : dout_r <= 12'hA2B;
			12'h74E : dout_r <= 12'hA28;
			12'h74F : dout_r <= 12'hA24;
			12'h750 : dout_r <= 12'hA21;
			12'h751 : dout_r <= 12'hA1E;
			12'h752 : dout_r <= 12'hA1B;
			12'h753 : dout_r <= 12'hA18;
			12'h754 : dout_r <= 12'hA15;
			12'h755 : dout_r <= 12'hA12;
			12'h756 : dout_r <= 12'hA0F;
			12'h757 : dout_r <= 12'hA0C;
			12'h758 : dout_r <= 12'hA09;
			12'h759 : dout_r <= 12'hA06;
			12'h75A : dout_r <= 12'hA03;
			12'h75B : dout_r <= 12'hA00;
			12'h75C : dout_r <= 12'h9FD;
			12'h75D : dout_r <= 12'h9FA;
			12'h75E : dout_r <= 12'h9F7;
			12'h75F : dout_r <= 12'h9F4;
			12'h760 : dout_r <= 12'h9F1;
			12'h761 : dout_r <= 12'h9EE;
			12'h762 : dout_r <= 12'h9EB;
			12'h763 : dout_r <= 12'h9E8;
			12'h764 : dout_r <= 12'h9E5;
			12'h765 : dout_r <= 12'h9E2;
			12'h766 : dout_r <= 12'h9DF;
			12'h767 : dout_r <= 12'h9DC;
			12'h768 : dout_r <= 12'h9D8;
			12'h769 : dout_r <= 12'h9D5;
			12'h76A : dout_r <= 12'h9D2;
			12'h76B : dout_r <= 12'h9CF;
			12'h76C : dout_r <= 12'h9CC;
			12'h76D : dout_r <= 12'h9C9;
			12'h76E : dout_r <= 12'h9C6;
			12'h76F : dout_r <= 12'h9C3;
			12'h770 : dout_r <= 12'h9C0;
			12'h771 : dout_r <= 12'h9BD;
			12'h772 : dout_r <= 12'h9BA;
			12'h773 : dout_r <= 12'h9B7;
			12'h774 : dout_r <= 12'h9B4;
			12'h775 : dout_r <= 12'h9B1;
			12'h776 : dout_r <= 12'h9AE;
			12'h777 : dout_r <= 12'h9AB;
			12'h778 : dout_r <= 12'h9A7;
			12'h779 : dout_r <= 12'h9A4;
			12'h77A : dout_r <= 12'h9A1;
			12'h77B : dout_r <= 12'h99E;
			12'h77C : dout_r <= 12'h99B;
			12'h77D : dout_r <= 12'h998;
			12'h77E : dout_r <= 12'h995;
			12'h77F : dout_r <= 12'h992;
			12'h780 : dout_r <= 12'h98F;
			12'h781 : dout_r <= 12'h98C;
			12'h782 : dout_r <= 12'h989;
			12'h783 : dout_r <= 12'h986;
			12'h784 : dout_r <= 12'h983;
			12'h785 : dout_r <= 12'h97F;
			12'h786 : dout_r <= 12'h97C;
			12'h787 : dout_r <= 12'h979;
			12'h788 : dout_r <= 12'h976;
			12'h789 : dout_r <= 12'h973;
			12'h78A : dout_r <= 12'h970;
			12'h78B : dout_r <= 12'h96D;
			12'h78C : dout_r <= 12'h96A;
			12'h78D : dout_r <= 12'h967;
			12'h78E : dout_r <= 12'h964;
			12'h78F : dout_r <= 12'h961;
			12'h790 : dout_r <= 12'h95D;
			12'h791 : dout_r <= 12'h95A;
			12'h792 : dout_r <= 12'h957;
			12'h793 : dout_r <= 12'h954;
			12'h794 : dout_r <= 12'h951;
			12'h795 : dout_r <= 12'h94E;
			12'h796 : dout_r <= 12'h94B;
			12'h797 : dout_r <= 12'h948;
			12'h798 : dout_r <= 12'h945;
			12'h799 : dout_r <= 12'h942;
			12'h79A : dout_r <= 12'h93E;
			12'h79B : dout_r <= 12'h93B;
			12'h79C : dout_r <= 12'h938;
			12'h79D : dout_r <= 12'h935;
			12'h79E : dout_r <= 12'h932;
			12'h79F : dout_r <= 12'h92F;
			12'h7A0 : dout_r <= 12'h92C;
			12'h7A1 : dout_r <= 12'h929;
			12'h7A2 : dout_r <= 12'h926;
			12'h7A3 : dout_r <= 12'h923;
			12'h7A4 : dout_r <= 12'h91F;
			12'h7A5 : dout_r <= 12'h91C;
			12'h7A6 : dout_r <= 12'h919;
			12'h7A7 : dout_r <= 12'h916;
			12'h7A8 : dout_r <= 12'h913;
			12'h7A9 : dout_r <= 12'h910;
			12'h7AA : dout_r <= 12'h90D;
			12'h7AB : dout_r <= 12'h90A;
			12'h7AC : dout_r <= 12'h907;
			12'h7AD : dout_r <= 12'h903;
			12'h7AE : dout_r <= 12'h900;
			12'h7AF : dout_r <= 12'h8FD;
			12'h7B0 : dout_r <= 12'h8FA;
			12'h7B1 : dout_r <= 12'h8F7;
			12'h7B2 : dout_r <= 12'h8F4;
			12'h7B3 : dout_r <= 12'h8F1;
			12'h7B4 : dout_r <= 12'h8EE;
			12'h7B5 : dout_r <= 12'h8EA;
			12'h7B6 : dout_r <= 12'h8E7;
			12'h7B7 : dout_r <= 12'h8E4;
			12'h7B8 : dout_r <= 12'h8E1;
			12'h7B9 : dout_r <= 12'h8DE;
			12'h7BA : dout_r <= 12'h8DB;
			12'h7BB : dout_r <= 12'h8D8;
			12'h7BC : dout_r <= 12'h8D5;
			12'h7BD : dout_r <= 12'h8D2;
			12'h7BE : dout_r <= 12'h8CE;
			12'h7BF : dout_r <= 12'h8CB;
			12'h7C0 : dout_r <= 12'h8C8;
			12'h7C1 : dout_r <= 12'h8C5;
			12'h7C2 : dout_r <= 12'h8C2;
			12'h7C3 : dout_r <= 12'h8BF;
			12'h7C4 : dout_r <= 12'h8BC;
			12'h7C5 : dout_r <= 12'h8B9;
			12'h7C6 : dout_r <= 12'h8B5;
			12'h7C7 : dout_r <= 12'h8B2;
			12'h7C8 : dout_r <= 12'h8AF;
			12'h7C9 : dout_r <= 12'h8AC;
			12'h7CA : dout_r <= 12'h8A9;
			12'h7CB : dout_r <= 12'h8A6;
			12'h7CC : dout_r <= 12'h8A3;
			12'h7CD : dout_r <= 12'h89F;
			12'h7CE : dout_r <= 12'h89C;
			12'h7CF : dout_r <= 12'h899;
			12'h7D0 : dout_r <= 12'h896;
			12'h7D1 : dout_r <= 12'h893;
			12'h7D2 : dout_r <= 12'h890;
			12'h7D3 : dout_r <= 12'h88D;
			12'h7D4 : dout_r <= 12'h88A;
			12'h7D5 : dout_r <= 12'h886;
			12'h7D6 : dout_r <= 12'h883;
			12'h7D7 : dout_r <= 12'h880;
			12'h7D8 : dout_r <= 12'h87D;
			12'h7D9 : dout_r <= 12'h87A;
			12'h7DA : dout_r <= 12'h877;
			12'h7DB : dout_r <= 12'h874;
			12'h7DC : dout_r <= 12'h870;
			12'h7DD : dout_r <= 12'h86D;
			12'h7DE : dout_r <= 12'h86A;
			12'h7DF : dout_r <= 12'h867;
			12'h7E0 : dout_r <= 12'h864;
			12'h7E1 : dout_r <= 12'h861;
			12'h7E2 : dout_r <= 12'h85E;
			12'h7E3 : dout_r <= 12'h85B;
			12'h7E4 : dout_r <= 12'h857;
			12'h7E5 : dout_r <= 12'h854;
			12'h7E6 : dout_r <= 12'h851;
			12'h7E7 : dout_r <= 12'h84E;
			12'h7E8 : dout_r <= 12'h84B;
			12'h7E9 : dout_r <= 12'h848;
			12'h7EA : dout_r <= 12'h845;
			12'h7EB : dout_r <= 12'h841;
			12'h7EC : dout_r <= 12'h83E;
			12'h7ED : dout_r <= 12'h83B;
			12'h7EE : dout_r <= 12'h838;
			12'h7EF : dout_r <= 12'h835;
			12'h7F0 : dout_r <= 12'h832;
			12'h7F1 : dout_r <= 12'h82F;
			12'h7F2 : dout_r <= 12'h82B;
			12'h7F3 : dout_r <= 12'h828;
			12'h7F4 : dout_r <= 12'h825;
			12'h7F5 : dout_r <= 12'h822;
			12'h7F6 : dout_r <= 12'h81F;
			12'h7F7 : dout_r <= 12'h81C;
			12'h7F8 : dout_r <= 12'h819;
			12'h7F9 : dout_r <= 12'h815;
			12'h7FA : dout_r <= 12'h812;
			12'h7FB : dout_r <= 12'h80F;
			12'h7FC : dout_r <= 12'h80C;
			12'h7FD : dout_r <= 12'h809;
			12'h7FE : dout_r <= 12'h806;
			12'h7FF : dout_r <= 12'h803;
			12'h800 : dout_r <= 12'h800;
			12'h801 : dout_r <= 12'h7FC;
			12'h802 : dout_r <= 12'h7F9;
			12'h803 : dout_r <= 12'h7F6;
			12'h804 : dout_r <= 12'h7F3;
			12'h805 : dout_r <= 12'h7F0;
			12'h806 : dout_r <= 12'h7ED;
			12'h807 : dout_r <= 12'h7EA;
			12'h808 : dout_r <= 12'h7E6;
			12'h809 : dout_r <= 12'h7E3;
			12'h80A : dout_r <= 12'h7E0;
			12'h80B : dout_r <= 12'h7DD;
			12'h80C : dout_r <= 12'h7DA;
			12'h80D : dout_r <= 12'h7D7;
			12'h80E : dout_r <= 12'h7D4;
			12'h80F : dout_r <= 12'h7D0;
			12'h810 : dout_r <= 12'h7CD;
			12'h811 : dout_r <= 12'h7CA;
			12'h812 : dout_r <= 12'h7C7;
			12'h813 : dout_r <= 12'h7C4;
			12'h814 : dout_r <= 12'h7C1;
			12'h815 : dout_r <= 12'h7BE;
			12'h816 : dout_r <= 12'h7BA;
			12'h817 : dout_r <= 12'h7B7;
			12'h818 : dout_r <= 12'h7B4;
			12'h819 : dout_r <= 12'h7B1;
			12'h81A : dout_r <= 12'h7AE;
			12'h81B : dout_r <= 12'h7AB;
			12'h81C : dout_r <= 12'h7A8;
			12'h81D : dout_r <= 12'h7A4;
			12'h81E : dout_r <= 12'h7A1;
			12'h81F : dout_r <= 12'h79E;
			12'h820 : dout_r <= 12'h79B;
			12'h821 : dout_r <= 12'h798;
			12'h822 : dout_r <= 12'h795;
			12'h823 : dout_r <= 12'h792;
			12'h824 : dout_r <= 12'h78F;
			12'h825 : dout_r <= 12'h78B;
			12'h826 : dout_r <= 12'h788;
			12'h827 : dout_r <= 12'h785;
			12'h828 : dout_r <= 12'h782;
			12'h829 : dout_r <= 12'h77F;
			12'h82A : dout_r <= 12'h77C;
			12'h82B : dout_r <= 12'h779;
			12'h82C : dout_r <= 12'h775;
			12'h82D : dout_r <= 12'h772;
			12'h82E : dout_r <= 12'h76F;
			12'h82F : dout_r <= 12'h76C;
			12'h830 : dout_r <= 12'h769;
			12'h831 : dout_r <= 12'h766;
			12'h832 : dout_r <= 12'h763;
			12'h833 : dout_r <= 12'h760;
			12'h834 : dout_r <= 12'h75C;
			12'h835 : dout_r <= 12'h759;
			12'h836 : dout_r <= 12'h756;
			12'h837 : dout_r <= 12'h753;
			12'h838 : dout_r <= 12'h750;
			12'h839 : dout_r <= 12'h74D;
			12'h83A : dout_r <= 12'h74A;
			12'h83B : dout_r <= 12'h746;
			12'h83C : dout_r <= 12'h743;
			12'h83D : dout_r <= 12'h740;
			12'h83E : dout_r <= 12'h73D;
			12'h83F : dout_r <= 12'h73A;
			12'h840 : dout_r <= 12'h737;
			12'h841 : dout_r <= 12'h734;
			12'h842 : dout_r <= 12'h731;
			12'h843 : dout_r <= 12'h72D;
			12'h844 : dout_r <= 12'h72A;
			12'h845 : dout_r <= 12'h727;
			12'h846 : dout_r <= 12'h724;
			12'h847 : dout_r <= 12'h721;
			12'h848 : dout_r <= 12'h71E;
			12'h849 : dout_r <= 12'h71B;
			12'h84A : dout_r <= 12'h718;
			12'h84B : dout_r <= 12'h715;
			12'h84C : dout_r <= 12'h711;
			12'h84D : dout_r <= 12'h70E;
			12'h84E : dout_r <= 12'h70B;
			12'h84F : dout_r <= 12'h708;
			12'h850 : dout_r <= 12'h705;
			12'h851 : dout_r <= 12'h702;
			12'h852 : dout_r <= 12'h6FF;
			12'h853 : dout_r <= 12'h6FC;
			12'h854 : dout_r <= 12'h6F8;
			12'h855 : dout_r <= 12'h6F5;
			12'h856 : dout_r <= 12'h6F2;
			12'h857 : dout_r <= 12'h6EF;
			12'h858 : dout_r <= 12'h6EC;
			12'h859 : dout_r <= 12'h6E9;
			12'h85A : dout_r <= 12'h6E6;
			12'h85B : dout_r <= 12'h6E3;
			12'h85C : dout_r <= 12'h6E0;
			12'h85D : dout_r <= 12'h6DC;
			12'h85E : dout_r <= 12'h6D9;
			12'h85F : dout_r <= 12'h6D6;
			12'h860 : dout_r <= 12'h6D3;
			12'h861 : dout_r <= 12'h6D0;
			12'h862 : dout_r <= 12'h6CD;
			12'h863 : dout_r <= 12'h6CA;
			12'h864 : dout_r <= 12'h6C7;
			12'h865 : dout_r <= 12'h6C4;
			12'h866 : dout_r <= 12'h6C1;
			12'h867 : dout_r <= 12'h6BD;
			12'h868 : dout_r <= 12'h6BA;
			12'h869 : dout_r <= 12'h6B7;
			12'h86A : dout_r <= 12'h6B4;
			12'h86B : dout_r <= 12'h6B1;
			12'h86C : dout_r <= 12'h6AE;
			12'h86D : dout_r <= 12'h6AB;
			12'h86E : dout_r <= 12'h6A8;
			12'h86F : dout_r <= 12'h6A5;
			12'h870 : dout_r <= 12'h6A2;
			12'h871 : dout_r <= 12'h69E;
			12'h872 : dout_r <= 12'h69B;
			12'h873 : dout_r <= 12'h698;
			12'h874 : dout_r <= 12'h695;
			12'h875 : dout_r <= 12'h692;
			12'h876 : dout_r <= 12'h68F;
			12'h877 : dout_r <= 12'h68C;
			12'h878 : dout_r <= 12'h689;
			12'h879 : dout_r <= 12'h686;
			12'h87A : dout_r <= 12'h683;
			12'h87B : dout_r <= 12'h680;
			12'h87C : dout_r <= 12'h67C;
			12'h87D : dout_r <= 12'h679;
			12'h87E : dout_r <= 12'h676;
			12'h87F : dout_r <= 12'h673;
			12'h880 : dout_r <= 12'h670;
			12'h881 : dout_r <= 12'h66D;
			12'h882 : dout_r <= 12'h66A;
			12'h883 : dout_r <= 12'h667;
			12'h884 : dout_r <= 12'h664;
			12'h885 : dout_r <= 12'h661;
			12'h886 : dout_r <= 12'h65E;
			12'h887 : dout_r <= 12'h65B;
			12'h888 : dout_r <= 12'h658;
			12'h889 : dout_r <= 12'h654;
			12'h88A : dout_r <= 12'h651;
			12'h88B : dout_r <= 12'h64E;
			12'h88C : dout_r <= 12'h64B;
			12'h88D : dout_r <= 12'h648;
			12'h88E : dout_r <= 12'h645;
			12'h88F : dout_r <= 12'h642;
			12'h890 : dout_r <= 12'h63F;
			12'h891 : dout_r <= 12'h63C;
			12'h892 : dout_r <= 12'h639;
			12'h893 : dout_r <= 12'h636;
			12'h894 : dout_r <= 12'h633;
			12'h895 : dout_r <= 12'h630;
			12'h896 : dout_r <= 12'h62D;
			12'h897 : dout_r <= 12'h62A;
			12'h898 : dout_r <= 12'h627;
			12'h899 : dout_r <= 12'h623;
			12'h89A : dout_r <= 12'h620;
			12'h89B : dout_r <= 12'h61D;
			12'h89C : dout_r <= 12'h61A;
			12'h89D : dout_r <= 12'h617;
			12'h89E : dout_r <= 12'h614;
			12'h89F : dout_r <= 12'h611;
			12'h8A0 : dout_r <= 12'h60E;
			12'h8A1 : dout_r <= 12'h60B;
			12'h8A2 : dout_r <= 12'h608;
			12'h8A3 : dout_r <= 12'h605;
			12'h8A4 : dout_r <= 12'h602;
			12'h8A5 : dout_r <= 12'h5FF;
			12'h8A6 : dout_r <= 12'h5FC;
			12'h8A7 : dout_r <= 12'h5F9;
			12'h8A8 : dout_r <= 12'h5F6;
			12'h8A9 : dout_r <= 12'h5F3;
			12'h8AA : dout_r <= 12'h5F0;
			12'h8AB : dout_r <= 12'h5ED;
			12'h8AC : dout_r <= 12'h5EA;
			12'h8AD : dout_r <= 12'h5E7;
			12'h8AE : dout_r <= 12'h5E4;
			12'h8AF : dout_r <= 12'h5E1;
			12'h8B0 : dout_r <= 12'h5DE;
			12'h8B1 : dout_r <= 12'h5DB;
			12'h8B2 : dout_r <= 12'h5D7;
			12'h8B3 : dout_r <= 12'h5D4;
			12'h8B4 : dout_r <= 12'h5D1;
			12'h8B5 : dout_r <= 12'h5CE;
			12'h8B6 : dout_r <= 12'h5CB;
			12'h8B7 : dout_r <= 12'h5C8;
			12'h8B8 : dout_r <= 12'h5C5;
			12'h8B9 : dout_r <= 12'h5C2;
			12'h8BA : dout_r <= 12'h5BF;
			12'h8BB : dout_r <= 12'h5BC;
			12'h8BC : dout_r <= 12'h5B9;
			12'h8BD : dout_r <= 12'h5B6;
			12'h8BE : dout_r <= 12'h5B3;
			12'h8BF : dout_r <= 12'h5B0;
			12'h8C0 : dout_r <= 12'h5AD;
			12'h8C1 : dout_r <= 12'h5AA;
			12'h8C2 : dout_r <= 12'h5A7;
			12'h8C3 : dout_r <= 12'h5A4;
			12'h8C4 : dout_r <= 12'h5A1;
			12'h8C5 : dout_r <= 12'h59E;
			12'h8C6 : dout_r <= 12'h59B;
			12'h8C7 : dout_r <= 12'h598;
			12'h8C8 : dout_r <= 12'h595;
			12'h8C9 : dout_r <= 12'h592;
			12'h8CA : dout_r <= 12'h58F;
			12'h8CB : dout_r <= 12'h58C;
			12'h8CC : dout_r <= 12'h589;
			12'h8CD : dout_r <= 12'h586;
			12'h8CE : dout_r <= 12'h583;
			12'h8CF : dout_r <= 12'h580;
			12'h8D0 : dout_r <= 12'h57D;
			12'h8D1 : dout_r <= 12'h57A;
			12'h8D2 : dout_r <= 12'h577;
			12'h8D3 : dout_r <= 12'h574;
			12'h8D4 : dout_r <= 12'h571;
			12'h8D5 : dout_r <= 12'h56F;
			12'h8D6 : dout_r <= 12'h56C;
			12'h8D7 : dout_r <= 12'h569;
			12'h8D8 : dout_r <= 12'h566;
			12'h8D9 : dout_r <= 12'h563;
			12'h8DA : dout_r <= 12'h560;
			12'h8DB : dout_r <= 12'h55D;
			12'h8DC : dout_r <= 12'h55A;
			12'h8DD : dout_r <= 12'h557;
			12'h8DE : dout_r <= 12'h554;
			12'h8DF : dout_r <= 12'h551;
			12'h8E0 : dout_r <= 12'h54E;
			12'h8E1 : dout_r <= 12'h54B;
			12'h8E2 : dout_r <= 12'h548;
			12'h8E3 : dout_r <= 12'h545;
			12'h8E4 : dout_r <= 12'h542;
			12'h8E5 : dout_r <= 12'h53F;
			12'h8E6 : dout_r <= 12'h53C;
			12'h8E7 : dout_r <= 12'h539;
			12'h8E8 : dout_r <= 12'h536;
			12'h8E9 : dout_r <= 12'h533;
			12'h8EA : dout_r <= 12'h530;
			12'h8EB : dout_r <= 12'h52D;
			12'h8EC : dout_r <= 12'h52B;
			12'h8ED : dout_r <= 12'h528;
			12'h8EE : dout_r <= 12'h525;
			12'h8EF : dout_r <= 12'h522;
			12'h8F0 : dout_r <= 12'h51F;
			12'h8F1 : dout_r <= 12'h51C;
			12'h8F2 : dout_r <= 12'h519;
			12'h8F3 : dout_r <= 12'h516;
			12'h8F4 : dout_r <= 12'h513;
			12'h8F5 : dout_r <= 12'h510;
			12'h8F6 : dout_r <= 12'h50D;
			12'h8F7 : dout_r <= 12'h50A;
			12'h8F8 : dout_r <= 12'h507;
			12'h8F9 : dout_r <= 12'h504;
			12'h8FA : dout_r <= 12'h502;
			12'h8FB : dout_r <= 12'h4FF;
			12'h8FC : dout_r <= 12'h4FC;
			12'h8FD : dout_r <= 12'h4F9;
			12'h8FE : dout_r <= 12'h4F6;
			12'h8FF : dout_r <= 12'h4F3;
			12'h900 : dout_r <= 12'h4F0;
			12'h901 : dout_r <= 12'h4ED;
			12'h902 : dout_r <= 12'h4EA;
			12'h903 : dout_r <= 12'h4E7;
			12'h904 : dout_r <= 12'h4E5;
			12'h905 : dout_r <= 12'h4E2;
			12'h906 : dout_r <= 12'h4DF;
			12'h907 : dout_r <= 12'h4DC;
			12'h908 : dout_r <= 12'h4D9;
			12'h909 : dout_r <= 12'h4D6;
			12'h90A : dout_r <= 12'h4D3;
			12'h90B : dout_r <= 12'h4D0;
			12'h90C : dout_r <= 12'h4CD;
			12'h90D : dout_r <= 12'h4CB;
			12'h90E : dout_r <= 12'h4C8;
			12'h90F : dout_r <= 12'h4C5;
			12'h910 : dout_r <= 12'h4C2;
			12'h911 : dout_r <= 12'h4BF;
			12'h912 : dout_r <= 12'h4BC;
			12'h913 : dout_r <= 12'h4B9;
			12'h914 : dout_r <= 12'h4B7;
			12'h915 : dout_r <= 12'h4B4;
			12'h916 : dout_r <= 12'h4B1;
			12'h917 : dout_r <= 12'h4AE;
			12'h918 : dout_r <= 12'h4AB;
			12'h919 : dout_r <= 12'h4A8;
			12'h91A : dout_r <= 12'h4A5;
			12'h91B : dout_r <= 12'h4A3;
			12'h91C : dout_r <= 12'h4A0;
			12'h91D : dout_r <= 12'h49D;
			12'h91E : dout_r <= 12'h49A;
			12'h91F : dout_r <= 12'h497;
			12'h920 : dout_r <= 12'h494;
			12'h921 : dout_r <= 12'h491;
			12'h922 : dout_r <= 12'h48F;
			12'h923 : dout_r <= 12'h48C;
			12'h924 : dout_r <= 12'h489;
			12'h925 : dout_r <= 12'h486;
			12'h926 : dout_r <= 12'h483;
			12'h927 : dout_r <= 12'h480;
			12'h928 : dout_r <= 12'h47E;
			12'h929 : dout_r <= 12'h47B;
			12'h92A : dout_r <= 12'h478;
			12'h92B : dout_r <= 12'h475;
			12'h92C : dout_r <= 12'h472;
			12'h92D : dout_r <= 12'h470;
			12'h92E : dout_r <= 12'h46D;
			12'h92F : dout_r <= 12'h46A;
			12'h930 : dout_r <= 12'h467;
			12'h931 : dout_r <= 12'h464;
			12'h932 : dout_r <= 12'h462;
			12'h933 : dout_r <= 12'h45F;
			12'h934 : dout_r <= 12'h45C;
			12'h935 : dout_r <= 12'h459;
			12'h936 : dout_r <= 12'h456;
			12'h937 : dout_r <= 12'h454;
			12'h938 : dout_r <= 12'h451;
			12'h939 : dout_r <= 12'h44E;
			12'h93A : dout_r <= 12'h44B;
			12'h93B : dout_r <= 12'h448;
			12'h93C : dout_r <= 12'h446;
			12'h93D : dout_r <= 12'h443;
			12'h93E : dout_r <= 12'h440;
			12'h93F : dout_r <= 12'h43D;
			12'h940 : dout_r <= 12'h43B;
			12'h941 : dout_r <= 12'h438;
			12'h942 : dout_r <= 12'h435;
			12'h943 : dout_r <= 12'h432;
			12'h944 : dout_r <= 12'h42F;
			12'h945 : dout_r <= 12'h42D;
			12'h946 : dout_r <= 12'h42A;
			12'h947 : dout_r <= 12'h427;
			12'h948 : dout_r <= 12'h424;
			12'h949 : dout_r <= 12'h422;
			12'h94A : dout_r <= 12'h41F;
			12'h94B : dout_r <= 12'h41C;
			12'h94C : dout_r <= 12'h419;
			12'h94D : dout_r <= 12'h417;
			12'h94E : dout_r <= 12'h414;
			12'h94F : dout_r <= 12'h411;
			12'h950 : dout_r <= 12'h40F;
			12'h951 : dout_r <= 12'h40C;
			12'h952 : dout_r <= 12'h409;
			12'h953 : dout_r <= 12'h406;
			12'h954 : dout_r <= 12'h404;
			12'h955 : dout_r <= 12'h401;
			12'h956 : dout_r <= 12'h3FE;
			12'h957 : dout_r <= 12'h3FB;
			12'h958 : dout_r <= 12'h3F9;
			12'h959 : dout_r <= 12'h3F6;
			12'h95A : dout_r <= 12'h3F3;
			12'h95B : dout_r <= 12'h3F1;
			12'h95C : dout_r <= 12'h3EE;
			12'h95D : dout_r <= 12'h3EB;
			12'h95E : dout_r <= 12'h3E9;
			12'h95F : dout_r <= 12'h3E6;
			12'h960 : dout_r <= 12'h3E3;
			12'h961 : dout_r <= 12'h3E0;
			12'h962 : dout_r <= 12'h3DE;
			12'h963 : dout_r <= 12'h3DB;
			12'h964 : dout_r <= 12'h3D8;
			12'h965 : dout_r <= 12'h3D6;
			12'h966 : dout_r <= 12'h3D3;
			12'h967 : dout_r <= 12'h3D0;
			12'h968 : dout_r <= 12'h3CE;
			12'h969 : dout_r <= 12'h3CB;
			12'h96A : dout_r <= 12'h3C8;
			12'h96B : dout_r <= 12'h3C6;
			12'h96C : dout_r <= 12'h3C3;
			12'h96D : dout_r <= 12'h3C0;
			12'h96E : dout_r <= 12'h3BE;
			12'h96F : dout_r <= 12'h3BB;
			12'h970 : dout_r <= 12'h3B8;
			12'h971 : dout_r <= 12'h3B6;
			12'h972 : dout_r <= 12'h3B3;
			12'h973 : dout_r <= 12'h3B0;
			12'h974 : dout_r <= 12'h3AE;
			12'h975 : dout_r <= 12'h3AB;
			12'h976 : dout_r <= 12'h3A8;
			12'h977 : dout_r <= 12'h3A6;
			12'h978 : dout_r <= 12'h3A3;
			12'h979 : dout_r <= 12'h3A1;
			12'h97A : dout_r <= 12'h39E;
			12'h97B : dout_r <= 12'h39B;
			12'h97C : dout_r <= 12'h399;
			12'h97D : dout_r <= 12'h396;
			12'h97E : dout_r <= 12'h393;
			12'h97F : dout_r <= 12'h391;
			12'h980 : dout_r <= 12'h38E;
			12'h981 : dout_r <= 12'h38C;
			12'h982 : dout_r <= 12'h389;
			12'h983 : dout_r <= 12'h386;
			12'h984 : dout_r <= 12'h384;
			12'h985 : dout_r <= 12'h381;
			12'h986 : dout_r <= 12'h37F;
			12'h987 : dout_r <= 12'h37C;
			12'h988 : dout_r <= 12'h379;
			12'h989 : dout_r <= 12'h377;
			12'h98A : dout_r <= 12'h374;
			12'h98B : dout_r <= 12'h372;
			12'h98C : dout_r <= 12'h36F;
			12'h98D : dout_r <= 12'h36D;
			12'h98E : dout_r <= 12'h36A;
			12'h98F : dout_r <= 12'h367;
			12'h990 : dout_r <= 12'h365;
			12'h991 : dout_r <= 12'h362;
			12'h992 : dout_r <= 12'h360;
			12'h993 : dout_r <= 12'h35D;
			12'h994 : dout_r <= 12'h35B;
			12'h995 : dout_r <= 12'h358;
			12'h996 : dout_r <= 12'h355;
			12'h997 : dout_r <= 12'h353;
			12'h998 : dout_r <= 12'h350;
			12'h999 : dout_r <= 12'h34E;
			12'h99A : dout_r <= 12'h34B;
			12'h99B : dout_r <= 12'h349;
			12'h99C : dout_r <= 12'h346;
			12'h99D : dout_r <= 12'h344;
			12'h99E : dout_r <= 12'h341;
			12'h99F : dout_r <= 12'h33F;
			12'h9A0 : dout_r <= 12'h33C;
			12'h9A1 : dout_r <= 12'h33A;
			12'h9A2 : dout_r <= 12'h337;
			12'h9A3 : dout_r <= 12'h335;
			12'h9A4 : dout_r <= 12'h332;
			12'h9A5 : dout_r <= 12'h330;
			12'h9A6 : dout_r <= 12'h32D;
			12'h9A7 : dout_r <= 12'h32B;
			12'h9A8 : dout_r <= 12'h328;
			12'h9A9 : dout_r <= 12'h326;
			12'h9AA : dout_r <= 12'h323;
			12'h9AB : dout_r <= 12'h321;
			12'h9AC : dout_r <= 12'h31E;
			12'h9AD : dout_r <= 12'h31C;
			12'h9AE : dout_r <= 12'h319;
			12'h9AF : dout_r <= 12'h317;
			12'h9B0 : dout_r <= 12'h314;
			12'h9B1 : dout_r <= 12'h312;
			12'h9B2 : dout_r <= 12'h30F;
			12'h9B3 : dout_r <= 12'h30D;
			12'h9B4 : dout_r <= 12'h30A;
			12'h9B5 : dout_r <= 12'h308;
			12'h9B6 : dout_r <= 12'h305;
			12'h9B7 : dout_r <= 12'h303;
			12'h9B8 : dout_r <= 12'h300;
			12'h9B9 : dout_r <= 12'h2FE;
			12'h9BA : dout_r <= 12'h2FC;
			12'h9BB : dout_r <= 12'h2F9;
			12'h9BC : dout_r <= 12'h2F7;
			12'h9BD : dout_r <= 12'h2F4;
			12'h9BE : dout_r <= 12'h2F2;
			12'h9BF : dout_r <= 12'h2EF;
			12'h9C0 : dout_r <= 12'h2ED;
			12'h9C1 : dout_r <= 12'h2EA;
			12'h9C2 : dout_r <= 12'h2E8;
			12'h9C3 : dout_r <= 12'h2E6;
			12'h9C4 : dout_r <= 12'h2E3;
			12'h9C5 : dout_r <= 12'h2E1;
			12'h9C6 : dout_r <= 12'h2DE;
			12'h9C7 : dout_r <= 12'h2DC;
			12'h9C8 : dout_r <= 12'h2DA;
			12'h9C9 : dout_r <= 12'h2D7;
			12'h9CA : dout_r <= 12'h2D5;
			12'h9CB : dout_r <= 12'h2D2;
			12'h9CC : dout_r <= 12'h2D0;
			12'h9CD : dout_r <= 12'h2CE;
			12'h9CE : dout_r <= 12'h2CB;
			12'h9CF : dout_r <= 12'h2C9;
			12'h9D0 : dout_r <= 12'h2C6;
			12'h9D1 : dout_r <= 12'h2C4;
			12'h9D2 : dout_r <= 12'h2C2;
			12'h9D3 : dout_r <= 12'h2BF;
			12'h9D4 : dout_r <= 12'h2BD;
			12'h9D5 : dout_r <= 12'h2BB;
			12'h9D6 : dout_r <= 12'h2B8;
			12'h9D7 : dout_r <= 12'h2B6;
			12'h9D8 : dout_r <= 12'h2B4;
			12'h9D9 : dout_r <= 12'h2B1;
			12'h9DA : dout_r <= 12'h2AF;
			12'h9DB : dout_r <= 12'h2AC;
			12'h9DC : dout_r <= 12'h2AA;
			12'h9DD : dout_r <= 12'h2A8;
			12'h9DE : dout_r <= 12'h2A5;
			12'h9DF : dout_r <= 12'h2A3;
			12'h9E0 : dout_r <= 12'h2A1;
			12'h9E1 : dout_r <= 12'h29E;
			12'h9E2 : dout_r <= 12'h29C;
			12'h9E3 : dout_r <= 12'h29A;
			12'h9E4 : dout_r <= 12'h298;
			12'h9E5 : dout_r <= 12'h295;
			12'h9E6 : dout_r <= 12'h293;
			12'h9E7 : dout_r <= 12'h291;
			12'h9E8 : dout_r <= 12'h28E;
			12'h9E9 : dout_r <= 12'h28C;
			12'h9EA : dout_r <= 12'h28A;
			12'h9EB : dout_r <= 12'h287;
			12'h9EC : dout_r <= 12'h285;
			12'h9ED : dout_r <= 12'h283;
			12'h9EE : dout_r <= 12'h281;
			12'h9EF : dout_r <= 12'h27E;
			12'h9F0 : dout_r <= 12'h27C;
			12'h9F1 : dout_r <= 12'h27A;
			12'h9F2 : dout_r <= 12'h277;
			12'h9F3 : dout_r <= 12'h275;
			12'h9F4 : dout_r <= 12'h273;
			12'h9F5 : dout_r <= 12'h271;
			12'h9F6 : dout_r <= 12'h26E;
			12'h9F7 : dout_r <= 12'h26C;
			12'h9F8 : dout_r <= 12'h26A;
			12'h9F9 : dout_r <= 12'h268;
			12'h9FA : dout_r <= 12'h265;
			12'h9FB : dout_r <= 12'h263;
			12'h9FC : dout_r <= 12'h261;
			12'h9FD : dout_r <= 12'h25F;
			12'h9FE : dout_r <= 12'h25C;
			12'h9FF : dout_r <= 12'h25A;
			12'hA00 : dout_r <= 12'h258;
			12'hA01 : dout_r <= 12'h256;
			12'hA02 : dout_r <= 12'h254;
			12'hA03 : dout_r <= 12'h251;
			12'hA04 : dout_r <= 12'h24F;
			12'hA05 : dout_r <= 12'h24D;
			12'hA06 : dout_r <= 12'h24B;
			12'hA07 : dout_r <= 12'h249;
			12'hA08 : dout_r <= 12'h246;
			12'hA09 : dout_r <= 12'h244;
			12'hA0A : dout_r <= 12'h242;
			12'hA0B : dout_r <= 12'h240;
			12'hA0C : dout_r <= 12'h23E;
			12'hA0D : dout_r <= 12'h23B;
			12'hA0E : dout_r <= 12'h239;
			12'hA0F : dout_r <= 12'h237;
			12'hA10 : dout_r <= 12'h235;
			12'hA11 : dout_r <= 12'h233;
			12'hA12 : dout_r <= 12'h231;
			12'hA13 : dout_r <= 12'h22E;
			12'hA14 : dout_r <= 12'h22C;
			12'hA15 : dout_r <= 12'h22A;
			12'hA16 : dout_r <= 12'h228;
			12'hA17 : dout_r <= 12'h226;
			12'hA18 : dout_r <= 12'h224;
			12'hA19 : dout_r <= 12'h222;
			12'hA1A : dout_r <= 12'h21F;
			12'hA1B : dout_r <= 12'h21D;
			12'hA1C : dout_r <= 12'h21B;
			12'hA1D : dout_r <= 12'h219;
			12'hA1E : dout_r <= 12'h217;
			12'hA1F : dout_r <= 12'h215;
			12'hA20 : dout_r <= 12'h213;
			12'hA21 : dout_r <= 12'h211;
			12'hA22 : dout_r <= 12'h20F;
			12'hA23 : dout_r <= 12'h20C;
			12'hA24 : dout_r <= 12'h20A;
			12'hA25 : dout_r <= 12'h208;
			12'hA26 : dout_r <= 12'h206;
			12'hA27 : dout_r <= 12'h204;
			12'hA28 : dout_r <= 12'h202;
			12'hA29 : dout_r <= 12'h200;
			12'hA2A : dout_r <= 12'h1FE;
			12'hA2B : dout_r <= 12'h1FC;
			12'hA2C : dout_r <= 12'h1FA;
			12'hA2D : dout_r <= 12'h1F8;
			12'hA2E : dout_r <= 12'h1F6;
			12'hA2F : dout_r <= 12'h1F4;
			12'hA30 : dout_r <= 12'h1F1;
			12'hA31 : dout_r <= 12'h1EF;
			12'hA32 : dout_r <= 12'h1ED;
			12'hA33 : dout_r <= 12'h1EB;
			12'hA34 : dout_r <= 12'h1E9;
			12'hA35 : dout_r <= 12'h1E7;
			12'hA36 : dout_r <= 12'h1E5;
			12'hA37 : dout_r <= 12'h1E3;
			12'hA38 : dout_r <= 12'h1E1;
			12'hA39 : dout_r <= 12'h1DF;
			12'hA3A : dout_r <= 12'h1DD;
			12'hA3B : dout_r <= 12'h1DB;
			12'hA3C : dout_r <= 12'h1D9;
			12'hA3D : dout_r <= 12'h1D7;
			12'hA3E : dout_r <= 12'h1D5;
			12'hA3F : dout_r <= 12'h1D3;
			12'hA40 : dout_r <= 12'h1D1;
			12'hA41 : dout_r <= 12'h1CF;
			12'hA42 : dout_r <= 12'h1CD;
			12'hA43 : dout_r <= 12'h1CB;
			12'hA44 : dout_r <= 12'h1C9;
			12'hA45 : dout_r <= 12'h1C7;
			12'hA46 : dout_r <= 12'h1C5;
			12'hA47 : dout_r <= 12'h1C3;
			12'hA48 : dout_r <= 12'h1C1;
			12'hA49 : dout_r <= 12'h1BF;
			12'hA4A : dout_r <= 12'h1BD;
			12'hA4B : dout_r <= 12'h1BB;
			12'hA4C : dout_r <= 12'h1BA;
			12'hA4D : dout_r <= 12'h1B8;
			12'hA4E : dout_r <= 12'h1B6;
			12'hA4F : dout_r <= 12'h1B4;
			12'hA50 : dout_r <= 12'h1B2;
			12'hA51 : dout_r <= 12'h1B0;
			12'hA52 : dout_r <= 12'h1AE;
			12'hA53 : dout_r <= 12'h1AC;
			12'hA54 : dout_r <= 12'h1AA;
			12'hA55 : dout_r <= 12'h1A8;
			12'hA56 : dout_r <= 12'h1A6;
			12'hA57 : dout_r <= 12'h1A4;
			12'hA58 : dout_r <= 12'h1A2;
			12'hA59 : dout_r <= 12'h1A1;
			12'hA5A : dout_r <= 12'h19F;
			12'hA5B : dout_r <= 12'h19D;
			12'hA5C : dout_r <= 12'h19B;
			12'hA5D : dout_r <= 12'h199;
			12'hA5E : dout_r <= 12'h197;
			12'hA5F : dout_r <= 12'h195;
			12'hA60 : dout_r <= 12'h193;
			12'hA61 : dout_r <= 12'h191;
			12'hA62 : dout_r <= 12'h190;
			12'hA63 : dout_r <= 12'h18E;
			12'hA64 : dout_r <= 12'h18C;
			12'hA65 : dout_r <= 12'h18A;
			12'hA66 : dout_r <= 12'h188;
			12'hA67 : dout_r <= 12'h186;
			12'hA68 : dout_r <= 12'h184;
			12'hA69 : dout_r <= 12'h183;
			12'hA6A : dout_r <= 12'h181;
			12'hA6B : dout_r <= 12'h17F;
			12'hA6C : dout_r <= 12'h17D;
			12'hA6D : dout_r <= 12'h17B;
			12'hA6E : dout_r <= 12'h17A;
			12'hA6F : dout_r <= 12'h178;
			12'hA70 : dout_r <= 12'h176;
			12'hA71 : dout_r <= 12'h174;
			12'hA72 : dout_r <= 12'h172;
			12'hA73 : dout_r <= 12'h170;
			12'hA74 : dout_r <= 12'h16F;
			12'hA75 : dout_r <= 12'h16D;
			12'hA76 : dout_r <= 12'h16B;
			12'hA77 : dout_r <= 12'h169;
			12'hA78 : dout_r <= 12'h168;
			12'hA79 : dout_r <= 12'h166;
			12'hA7A : dout_r <= 12'h164;
			12'hA7B : dout_r <= 12'h162;
			12'hA7C : dout_r <= 12'h160;
			12'hA7D : dout_r <= 12'h15F;
			12'hA7E : dout_r <= 12'h15D;
			12'hA7F : dout_r <= 12'h15B;
			12'hA80 : dout_r <= 12'h159;
			12'hA81 : dout_r <= 12'h158;
			12'hA82 : dout_r <= 12'h156;
			12'hA83 : dout_r <= 12'h154;
			12'hA84 : dout_r <= 12'h153;
			12'hA85 : dout_r <= 12'h151;
			12'hA86 : dout_r <= 12'h14F;
			12'hA87 : dout_r <= 12'h14D;
			12'hA88 : dout_r <= 12'h14C;
			12'hA89 : dout_r <= 12'h14A;
			12'hA8A : dout_r <= 12'h148;
			12'hA8B : dout_r <= 12'h147;
			12'hA8C : dout_r <= 12'h145;
			12'hA8D : dout_r <= 12'h143;
			12'hA8E : dout_r <= 12'h141;
			12'hA8F : dout_r <= 12'h140;
			12'hA90 : dout_r <= 12'h13E;
			12'hA91 : dout_r <= 12'h13C;
			12'hA92 : dout_r <= 12'h13B;
			12'hA93 : dout_r <= 12'h139;
			12'hA94 : dout_r <= 12'h137;
			12'hA95 : dout_r <= 12'h136;
			12'hA96 : dout_r <= 12'h134;
			12'hA97 : dout_r <= 12'h132;
			12'hA98 : dout_r <= 12'h131;
			12'hA99 : dout_r <= 12'h12F;
			12'hA9A : dout_r <= 12'h12D;
			12'hA9B : dout_r <= 12'h12C;
			12'hA9C : dout_r <= 12'h12A;
			12'hA9D : dout_r <= 12'h129;
			12'hA9E : dout_r <= 12'h127;
			12'hA9F : dout_r <= 12'h125;
			12'hAA0 : dout_r <= 12'h124;
			12'hAA1 : dout_r <= 12'h122;
			12'hAA2 : dout_r <= 12'h121;
			12'hAA3 : dout_r <= 12'h11F;
			12'hAA4 : dout_r <= 12'h11D;
			12'hAA5 : dout_r <= 12'h11C;
			12'hAA6 : dout_r <= 12'h11A;
			12'hAA7 : dout_r <= 12'h119;
			12'hAA8 : dout_r <= 12'h117;
			12'hAA9 : dout_r <= 12'h115;
			12'hAAA : dout_r <= 12'h114;
			12'hAAB : dout_r <= 12'h112;
			12'hAAC : dout_r <= 12'h111;
			12'hAAD : dout_r <= 12'h10F;
			12'hAAE : dout_r <= 12'h10E;
			12'hAAF : dout_r <= 12'h10C;
			12'hAB0 : dout_r <= 12'h10A;
			12'hAB1 : dout_r <= 12'h109;
			12'hAB2 : dout_r <= 12'h107;
			12'hAB3 : dout_r <= 12'h106;
			12'hAB4 : dout_r <= 12'h104;
			12'hAB5 : dout_r <= 12'h103;
			12'hAB6 : dout_r <= 12'h101;
			12'hAB7 : dout_r <= 12'h100;
			12'hAB8 : dout_r <= 12'h0FE;
			12'hAB9 : dout_r <= 12'h0FD;
			12'hABA : dout_r <= 12'h0FB;
			12'hABB : dout_r <= 12'h0FA;
			12'hABC : dout_r <= 12'h0F8;
			12'hABD : dout_r <= 12'h0F7;
			12'hABE : dout_r <= 12'h0F5;
			12'hABF : dout_r <= 12'h0F4;
			12'hAC0 : dout_r <= 12'h0F2;
			12'hAC1 : dout_r <= 12'h0F1;
			12'hAC2 : dout_r <= 12'h0EF;
			12'hAC3 : dout_r <= 12'h0EE;
			12'hAC4 : dout_r <= 12'h0EC;
			12'hAC5 : dout_r <= 12'h0EB;
			12'hAC6 : dout_r <= 12'h0E9;
			12'hAC7 : dout_r <= 12'h0E8;
			12'hAC8 : dout_r <= 12'h0E7;
			12'hAC9 : dout_r <= 12'h0E5;
			12'hACA : dout_r <= 12'h0E4;
			12'hACB : dout_r <= 12'h0E2;
			12'hACC : dout_r <= 12'h0E1;
			12'hACD : dout_r <= 12'h0DF;
			12'hACE : dout_r <= 12'h0DE;
			12'hACF : dout_r <= 12'h0DC;
			12'hAD0 : dout_r <= 12'h0DB;
			12'hAD1 : dout_r <= 12'h0DA;
			12'hAD2 : dout_r <= 12'h0D8;
			12'hAD3 : dout_r <= 12'h0D7;
			12'hAD4 : dout_r <= 12'h0D5;
			12'hAD5 : dout_r <= 12'h0D4;
			12'hAD6 : dout_r <= 12'h0D3;
			12'hAD7 : dout_r <= 12'h0D1;
			12'hAD8 : dout_r <= 12'h0D0;
			12'hAD9 : dout_r <= 12'h0CF;
			12'hADA : dout_r <= 12'h0CD;
			12'hADB : dout_r <= 12'h0CC;
			12'hADC : dout_r <= 12'h0CA;
			12'hADD : dout_r <= 12'h0C9;
			12'hADE : dout_r <= 12'h0C8;
			12'hADF : dout_r <= 12'h0C6;
			12'hAE0 : dout_r <= 12'h0C5;
			12'hAE1 : dout_r <= 12'h0C4;
			12'hAE2 : dout_r <= 12'h0C2;
			12'hAE3 : dout_r <= 12'h0C1;
			12'hAE4 : dout_r <= 12'h0C0;
			12'hAE5 : dout_r <= 12'h0BE;
			12'hAE6 : dout_r <= 12'h0BD;
			12'hAE7 : dout_r <= 12'h0BC;
			12'hAE8 : dout_r <= 12'h0BA;
			12'hAE9 : dout_r <= 12'h0B9;
			12'hAEA : dout_r <= 12'h0B8;
			12'hAEB : dout_r <= 12'h0B7;
			12'hAEC : dout_r <= 12'h0B5;
			12'hAED : dout_r <= 12'h0B4;
			12'hAEE : dout_r <= 12'h0B3;
			12'hAEF : dout_r <= 12'h0B1;
			12'hAF0 : dout_r <= 12'h0B0;
			12'hAF1 : dout_r <= 12'h0AF;
			12'hAF2 : dout_r <= 12'h0AE;
			12'hAF3 : dout_r <= 12'h0AC;
			12'hAF4 : dout_r <= 12'h0AB;
			12'hAF5 : dout_r <= 12'h0AA;
			12'hAF6 : dout_r <= 12'h0A9;
			12'hAF7 : dout_r <= 12'h0A7;
			12'hAF8 : dout_r <= 12'h0A6;
			12'hAF9 : dout_r <= 12'h0A5;
			12'hAFA : dout_r <= 12'h0A4;
			12'hAFB : dout_r <= 12'h0A2;
			12'hAFC : dout_r <= 12'h0A1;
			12'hAFD : dout_r <= 12'h0A0;
			12'hAFE : dout_r <= 12'h09F;
			12'hAFF : dout_r <= 12'h09E;
			12'hB00 : dout_r <= 12'h09C;
			12'hB01 : dout_r <= 12'h09B;
			12'hB02 : dout_r <= 12'h09A;
			12'hB03 : dout_r <= 12'h099;
			12'hB04 : dout_r <= 12'h098;
			12'hB05 : dout_r <= 12'h096;
			12'hB06 : dout_r <= 12'h095;
			12'hB07 : dout_r <= 12'h094;
			12'hB08 : dout_r <= 12'h093;
			12'hB09 : dout_r <= 12'h092;
			12'hB0A : dout_r <= 12'h091;
			12'hB0B : dout_r <= 12'h08F;
			12'hB0C : dout_r <= 12'h08E;
			12'hB0D : dout_r <= 12'h08D;
			12'hB0E : dout_r <= 12'h08C;
			12'hB0F : dout_r <= 12'h08B;
			12'hB10 : dout_r <= 12'h08A;
			12'hB11 : dout_r <= 12'h089;
			12'hB12 : dout_r <= 12'h087;
			12'hB13 : dout_r <= 12'h086;
			12'hB14 : dout_r <= 12'h085;
			12'hB15 : dout_r <= 12'h084;
			12'hB16 : dout_r <= 12'h083;
			12'hB17 : dout_r <= 12'h082;
			12'hB18 : dout_r <= 12'h081;
			12'hB19 : dout_r <= 12'h080;
			12'hB1A : dout_r <= 12'h07F;
			12'hB1B : dout_r <= 12'h07E;
			12'hB1C : dout_r <= 12'h07C;
			12'hB1D : dout_r <= 12'h07B;
			12'hB1E : dout_r <= 12'h07A;
			12'hB1F : dout_r <= 12'h079;
			12'hB20 : dout_r <= 12'h078;
			12'hB21 : dout_r <= 12'h077;
			12'hB22 : dout_r <= 12'h076;
			12'hB23 : dout_r <= 12'h075;
			12'hB24 : dout_r <= 12'h074;
			12'hB25 : dout_r <= 12'h073;
			12'hB26 : dout_r <= 12'h072;
			12'hB27 : dout_r <= 12'h071;
			12'hB28 : dout_r <= 12'h070;
			12'hB29 : dout_r <= 12'h06F;
			12'hB2A : dout_r <= 12'h06E;
			12'hB2B : dout_r <= 12'h06D;
			12'hB2C : dout_r <= 12'h06C;
			12'hB2D : dout_r <= 12'h06B;
			12'hB2E : dout_r <= 12'h06A;
			12'hB2F : dout_r <= 12'h069;
			12'hB30 : dout_r <= 12'h068;
			12'hB31 : dout_r <= 12'h067;
			12'hB32 : dout_r <= 12'h066;
			12'hB33 : dout_r <= 12'h065;
			12'hB34 : dout_r <= 12'h064;
			12'hB35 : dout_r <= 12'h063;
			12'hB36 : dout_r <= 12'h062;
			12'hB37 : dout_r <= 12'h061;
			12'hB38 : dout_r <= 12'h060;
			12'hB39 : dout_r <= 12'h05F;
			12'hB3A : dout_r <= 12'h05E;
			12'hB3B : dout_r <= 12'h05D;
			12'hB3C : dout_r <= 12'h05C;
			12'hB3D : dout_r <= 12'h05B;
			12'hB3E : dout_r <= 12'h05A;
			12'hB3F : dout_r <= 12'h05A;
			12'hB40 : dout_r <= 12'h059;
			12'hB41 : dout_r <= 12'h058;
			12'hB42 : dout_r <= 12'h057;
			12'hB43 : dout_r <= 12'h056;
			12'hB44 : dout_r <= 12'h055;
			12'hB45 : dout_r <= 12'h054;
			12'hB46 : dout_r <= 12'h053;
			12'hB47 : dout_r <= 12'h052;
			12'hB48 : dout_r <= 12'h051;
			12'hB49 : dout_r <= 12'h051;
			12'hB4A : dout_r <= 12'h050;
			12'hB4B : dout_r <= 12'h04F;
			12'hB4C : dout_r <= 12'h04E;
			12'hB4D : dout_r <= 12'h04D;
			12'hB4E : dout_r <= 12'h04C;
			12'hB4F : dout_r <= 12'h04B;
			12'hB50 : dout_r <= 12'h04B;
			12'hB51 : dout_r <= 12'h04A;
			12'hB52 : dout_r <= 12'h049;
			12'hB53 : dout_r <= 12'h048;
			12'hB54 : dout_r <= 12'h047;
			12'hB55 : dout_r <= 12'h047;
			12'hB56 : dout_r <= 12'h046;
			12'hB57 : dout_r <= 12'h045;
			12'hB58 : dout_r <= 12'h044;
			12'hB59 : dout_r <= 12'h043;
			12'hB5A : dout_r <= 12'h043;
			12'hB5B : dout_r <= 12'h042;
			12'hB5C : dout_r <= 12'h041;
			12'hB5D : dout_r <= 12'h040;
			12'hB5E : dout_r <= 12'h03F;
			12'hB5F : dout_r <= 12'h03F;
			12'hB60 : dout_r <= 12'h03E;
			12'hB61 : dout_r <= 12'h03D;
			12'hB62 : dout_r <= 12'h03C;
			12'hB63 : dout_r <= 12'h03C;
			12'hB64 : dout_r <= 12'h03B;
			12'hB65 : dout_r <= 12'h03A;
			12'hB66 : dout_r <= 12'h039;
			12'hB67 : dout_r <= 12'h039;
			12'hB68 : dout_r <= 12'h038;
			12'hB69 : dout_r <= 12'h037;
			12'hB6A : dout_r <= 12'h036;
			12'hB6B : dout_r <= 12'h036;
			12'hB6C : dout_r <= 12'h035;
			12'hB6D : dout_r <= 12'h034;
			12'hB6E : dout_r <= 12'h034;
			12'hB6F : dout_r <= 12'h033;
			12'hB70 : dout_r <= 12'h032;
			12'hB71 : dout_r <= 12'h032;
			12'hB72 : dout_r <= 12'h031;
			12'hB73 : dout_r <= 12'h030;
			12'hB74 : dout_r <= 12'h030;
			12'hB75 : dout_r <= 12'h02F;
			12'hB76 : dout_r <= 12'h02E;
			12'hB77 : dout_r <= 12'h02E;
			12'hB78 : dout_r <= 12'h02D;
			12'hB79 : dout_r <= 12'h02C;
			12'hB7A : dout_r <= 12'h02C;
			12'hB7B : dout_r <= 12'h02B;
			12'hB7C : dout_r <= 12'h02A;
			12'hB7D : dout_r <= 12'h02A;
			12'hB7E : dout_r <= 12'h029;
			12'hB7F : dout_r <= 12'h028;
			12'hB80 : dout_r <= 12'h028;
			12'hB81 : dout_r <= 12'h027;
			12'hB82 : dout_r <= 12'h027;
			12'hB83 : dout_r <= 12'h026;
			12'hB84 : dout_r <= 12'h025;
			12'hB85 : dout_r <= 12'h025;
			12'hB86 : dout_r <= 12'h024;
			12'hB87 : dout_r <= 12'h024;
			12'hB88 : dout_r <= 12'h023;
			12'hB89 : dout_r <= 12'h023;
			12'hB8A : dout_r <= 12'h022;
			12'hB8B : dout_r <= 12'h021;
			12'hB8C : dout_r <= 12'h021;
			12'hB8D : dout_r <= 12'h020;
			12'hB8E : dout_r <= 12'h020;
			12'hB8F : dout_r <= 12'h01F;
			12'hB90 : dout_r <= 12'h01F;
			12'hB91 : dout_r <= 12'h01E;
			12'hB92 : dout_r <= 12'h01E;
			12'hB93 : dout_r <= 12'h01D;
			12'hB94 : dout_r <= 12'h01D;
			12'hB95 : dout_r <= 12'h01C;
			12'hB96 : dout_r <= 12'h01C;
			12'hB97 : dout_r <= 12'h01B;
			12'hB98 : dout_r <= 12'h01A;
			12'hB99 : dout_r <= 12'h01A;
			12'hB9A : dout_r <= 12'h01A;
			12'hB9B : dout_r <= 12'h019;
			12'hB9C : dout_r <= 12'h019;
			12'hB9D : dout_r <= 12'h018;
			12'hB9E : dout_r <= 12'h018;
			12'hB9F : dout_r <= 12'h017;
			12'hBA0 : dout_r <= 12'h017;
			12'hBA1 : dout_r <= 12'h016;
			12'hBA2 : dout_r <= 12'h016;
			12'hBA3 : dout_r <= 12'h015;
			12'hBA4 : dout_r <= 12'h015;
			12'hBA5 : dout_r <= 12'h014;
			12'hBA6 : dout_r <= 12'h014;
			12'hBA7 : dout_r <= 12'h014;
			12'hBA8 : dout_r <= 12'h013;
			12'hBA9 : dout_r <= 12'h013;
			12'hBAA : dout_r <= 12'h012;
			12'hBAB : dout_r <= 12'h012;
			12'hBAC : dout_r <= 12'h011;
			12'hBAD : dout_r <= 12'h011;
			12'hBAE : dout_r <= 12'h011;
			12'hBAF : dout_r <= 12'h010;
			12'hBB0 : dout_r <= 12'h010;
			12'hBB1 : dout_r <= 12'h010;
			12'hBB2 : dout_r <= 12'h00F;
			12'hBB3 : dout_r <= 12'h00F;
			12'hBB4 : dout_r <= 12'h00E;
			12'hBB5 : dout_r <= 12'h00E;
			12'hBB6 : dout_r <= 12'h00E;
			12'hBB7 : dout_r <= 12'h00D;
			12'hBB8 : dout_r <= 12'h00D;
			12'hBB9 : dout_r <= 12'h00D;
			12'hBBA : dout_r <= 12'h00C;
			12'hBBB : dout_r <= 12'h00C;
			12'hBBC : dout_r <= 12'h00C;
			12'hBBD : dout_r <= 12'h00B;
			12'hBBE : dout_r <= 12'h00B;
			12'hBBF : dout_r <= 12'h00B;
			12'hBC0 : dout_r <= 12'h00A;
			12'hBC1 : dout_r <= 12'h00A;
			12'hBC2 : dout_r <= 12'h00A;
			12'hBC3 : dout_r <= 12'h009;
			12'hBC4 : dout_r <= 12'h009;
			12'hBC5 : dout_r <= 12'h009;
			12'hBC6 : dout_r <= 12'h009;
			12'hBC7 : dout_r <= 12'h008;
			12'hBC8 : dout_r <= 12'h008;
			12'hBC9 : dout_r <= 12'h008;
			12'hBCA : dout_r <= 12'h008;
			12'hBCB : dout_r <= 12'h007;
			12'hBCC : dout_r <= 12'h007;
			12'hBCD : dout_r <= 12'h007;
			12'hBCE : dout_r <= 12'h007;
			12'hBCF : dout_r <= 12'h006;
			12'hBD0 : dout_r <= 12'h006;
			12'hBD1 : dout_r <= 12'h006;
			12'hBD2 : dout_r <= 12'h006;
			12'hBD3 : dout_r <= 12'h005;
			12'hBD4 : dout_r <= 12'h005;
			12'hBD5 : dout_r <= 12'h005;
			12'hBD6 : dout_r <= 12'h005;
			12'hBD7 : dout_r <= 12'h005;
			12'hBD8 : dout_r <= 12'h004;
			12'hBD9 : dout_r <= 12'h004;
			12'hBDA : dout_r <= 12'h004;
			12'hBDB : dout_r <= 12'h004;
			12'hBDC : dout_r <= 12'h004;
			12'hBDD : dout_r <= 12'h003;
			12'hBDE : dout_r <= 12'h003;
			12'hBDF : dout_r <= 12'h003;
			12'hBE0 : dout_r <= 12'h003;
			12'hBE1 : dout_r <= 12'h003;
			12'hBE2 : dout_r <= 12'h003;
			12'hBE3 : dout_r <= 12'h003;
			12'hBE4 : dout_r <= 12'h002;
			12'hBE5 : dout_r <= 12'h002;
			12'hBE6 : dout_r <= 12'h002;
			12'hBE7 : dout_r <= 12'h002;
			12'hBE8 : dout_r <= 12'h002;
			12'hBE9 : dout_r <= 12'h002;
			12'hBEA : dout_r <= 12'h002;
			12'hBEB : dout_r <= 12'h002;
			12'hBEC : dout_r <= 12'h001;
			12'hBED : dout_r <= 12'h001;
			12'hBEE : dout_r <= 12'h001;
			12'hBEF : dout_r <= 12'h001;
			12'hBF0 : dout_r <= 12'h001;
			12'hBF1 : dout_r <= 12'h001;
			12'hBF2 : dout_r <= 12'h001;
			12'hBF3 : dout_r <= 12'h001;
			12'hBF4 : dout_r <= 12'h001;
			12'hBF5 : dout_r <= 12'h001;
			12'hBF6 : dout_r <= 12'h001;
			12'hBF7 : dout_r <= 12'h001;
			12'hBF8 : dout_r <= 12'h001;
			12'hBF9 : dout_r <= 12'h001;
			12'hBFA : dout_r <= 12'h001;
			12'hBFB : dout_r <= 12'h001;
			12'hBFC : dout_r <= 12'h001;
			12'hBFD : dout_r <= 12'h001;
			12'hBFE : dout_r <= 12'h001;
			12'hBFF : dout_r <= 12'h001;
			12'hC00 : dout_r <= 12'h000;
			12'hC01 : dout_r <= 12'h001;
			12'hC02 : dout_r <= 12'h001;
			12'hC03 : dout_r <= 12'h001;
			12'hC04 : dout_r <= 12'h001;
			12'hC05 : dout_r <= 12'h001;
			12'hC06 : dout_r <= 12'h001;
			12'hC07 : dout_r <= 12'h001;
			12'hC08 : dout_r <= 12'h001;
			12'hC09 : dout_r <= 12'h001;
			12'hC0A : dout_r <= 12'h001;
			12'hC0B : dout_r <= 12'h001;
			12'hC0C : dout_r <= 12'h001;
			12'hC0D : dout_r <= 12'h001;
			12'hC0E : dout_r <= 12'h001;
			12'hC0F : dout_r <= 12'h001;
			12'hC10 : dout_r <= 12'h001;
			12'hC11 : dout_r <= 12'h001;
			12'hC12 : dout_r <= 12'h001;
			12'hC13 : dout_r <= 12'h001;
			12'hC14 : dout_r <= 12'h001;
			12'hC15 : dout_r <= 12'h002;
			12'hC16 : dout_r <= 12'h002;
			12'hC17 : dout_r <= 12'h002;
			12'hC18 : dout_r <= 12'h002;
			12'hC19 : dout_r <= 12'h002;
			12'hC1A : dout_r <= 12'h002;
			12'hC1B : dout_r <= 12'h002;
			12'hC1C : dout_r <= 12'h002;
			12'hC1D : dout_r <= 12'h003;
			12'hC1E : dout_r <= 12'h003;
			12'hC1F : dout_r <= 12'h003;
			12'hC20 : dout_r <= 12'h003;
			12'hC21 : dout_r <= 12'h003;
			12'hC22 : dout_r <= 12'h003;
			12'hC23 : dout_r <= 12'h003;
			12'hC24 : dout_r <= 12'h004;
			12'hC25 : dout_r <= 12'h004;
			12'hC26 : dout_r <= 12'h004;
			12'hC27 : dout_r <= 12'h004;
			12'hC28 : dout_r <= 12'h004;
			12'hC29 : dout_r <= 12'h005;
			12'hC2A : dout_r <= 12'h005;
			12'hC2B : dout_r <= 12'h005;
			12'hC2C : dout_r <= 12'h005;
			12'hC2D : dout_r <= 12'h005;
			12'hC2E : dout_r <= 12'h006;
			12'hC2F : dout_r <= 12'h006;
			12'hC30 : dout_r <= 12'h006;
			12'hC31 : dout_r <= 12'h006;
			12'hC32 : dout_r <= 12'h007;
			12'hC33 : dout_r <= 12'h007;
			12'hC34 : dout_r <= 12'h007;
			12'hC35 : dout_r <= 12'h007;
			12'hC36 : dout_r <= 12'h008;
			12'hC37 : dout_r <= 12'h008;
			12'hC38 : dout_r <= 12'h008;
			12'hC39 : dout_r <= 12'h008;
			12'hC3A : dout_r <= 12'h009;
			12'hC3B : dout_r <= 12'h009;
			12'hC3C : dout_r <= 12'h009;
			12'hC3D : dout_r <= 12'h009;
			12'hC3E : dout_r <= 12'h00A;
			12'hC3F : dout_r <= 12'h00A;
			12'hC40 : dout_r <= 12'h00A;
			12'hC41 : dout_r <= 12'h00B;
			12'hC42 : dout_r <= 12'h00B;
			12'hC43 : dout_r <= 12'h00B;
			12'hC44 : dout_r <= 12'h00C;
			12'hC45 : dout_r <= 12'h00C;
			12'hC46 : dout_r <= 12'h00C;
			12'hC47 : dout_r <= 12'h00D;
			12'hC48 : dout_r <= 12'h00D;
			12'hC49 : dout_r <= 12'h00D;
			12'hC4A : dout_r <= 12'h00E;
			12'hC4B : dout_r <= 12'h00E;
			12'hC4C : dout_r <= 12'h00E;
			12'hC4D : dout_r <= 12'h00F;
			12'hC4E : dout_r <= 12'h00F;
			12'hC4F : dout_r <= 12'h010;
			12'hC50 : dout_r <= 12'h010;
			12'hC51 : dout_r <= 12'h010;
			12'hC52 : dout_r <= 12'h011;
			12'hC53 : dout_r <= 12'h011;
			12'hC54 : dout_r <= 12'h011;
			12'hC55 : dout_r <= 12'h012;
			12'hC56 : dout_r <= 12'h012;
			12'hC57 : dout_r <= 12'h013;
			12'hC58 : dout_r <= 12'h013;
			12'hC59 : dout_r <= 12'h014;
			12'hC5A : dout_r <= 12'h014;
			12'hC5B : dout_r <= 12'h014;
			12'hC5C : dout_r <= 12'h015;
			12'hC5D : dout_r <= 12'h015;
			12'hC5E : dout_r <= 12'h016;
			12'hC5F : dout_r <= 12'h016;
			12'hC60 : dout_r <= 12'h017;
			12'hC61 : dout_r <= 12'h017;
			12'hC62 : dout_r <= 12'h018;
			12'hC63 : dout_r <= 12'h018;
			12'hC64 : dout_r <= 12'h019;
			12'hC65 : dout_r <= 12'h019;
			12'hC66 : dout_r <= 12'h01A;
			12'hC67 : dout_r <= 12'h01A;
			12'hC68 : dout_r <= 12'h01A;
			12'hC69 : dout_r <= 12'h01B;
			12'hC6A : dout_r <= 12'h01C;
			12'hC6B : dout_r <= 12'h01C;
			12'hC6C : dout_r <= 12'h01D;
			12'hC6D : dout_r <= 12'h01D;
			12'hC6E : dout_r <= 12'h01E;
			12'hC6F : dout_r <= 12'h01E;
			12'hC70 : dout_r <= 12'h01F;
			12'hC71 : dout_r <= 12'h01F;
			12'hC72 : dout_r <= 12'h020;
			12'hC73 : dout_r <= 12'h020;
			12'hC74 : dout_r <= 12'h021;
			12'hC75 : dout_r <= 12'h021;
			12'hC76 : dout_r <= 12'h022;
			12'hC77 : dout_r <= 12'h023;
			12'hC78 : dout_r <= 12'h023;
			12'hC79 : dout_r <= 12'h024;
			12'hC7A : dout_r <= 12'h024;
			12'hC7B : dout_r <= 12'h025;
			12'hC7C : dout_r <= 12'h025;
			12'hC7D : dout_r <= 12'h026;
			12'hC7E : dout_r <= 12'h027;
			12'hC7F : dout_r <= 12'h027;
			12'hC80 : dout_r <= 12'h028;
			12'hC81 : dout_r <= 12'h028;
			12'hC82 : dout_r <= 12'h029;
			12'hC83 : dout_r <= 12'h02A;
			12'hC84 : dout_r <= 12'h02A;
			12'hC85 : dout_r <= 12'h02B;
			12'hC86 : dout_r <= 12'h02C;
			12'hC87 : dout_r <= 12'h02C;
			12'hC88 : dout_r <= 12'h02D;
			12'hC89 : dout_r <= 12'h02E;
			12'hC8A : dout_r <= 12'h02E;
			12'hC8B : dout_r <= 12'h02F;
			12'hC8C : dout_r <= 12'h030;
			12'hC8D : dout_r <= 12'h030;
			12'hC8E : dout_r <= 12'h031;
			12'hC8F : dout_r <= 12'h032;
			12'hC90 : dout_r <= 12'h032;
			12'hC91 : dout_r <= 12'h033;
			12'hC92 : dout_r <= 12'h034;
			12'hC93 : dout_r <= 12'h034;
			12'hC94 : dout_r <= 12'h035;
			12'hC95 : dout_r <= 12'h036;
			12'hC96 : dout_r <= 12'h036;
			12'hC97 : dout_r <= 12'h037;
			12'hC98 : dout_r <= 12'h038;
			12'hC99 : dout_r <= 12'h039;
			12'hC9A : dout_r <= 12'h039;
			12'hC9B : dout_r <= 12'h03A;
			12'hC9C : dout_r <= 12'h03B;
			12'hC9D : dout_r <= 12'h03C;
			12'hC9E : dout_r <= 12'h03C;
			12'hC9F : dout_r <= 12'h03D;
			12'hCA0 : dout_r <= 12'h03E;
			12'hCA1 : dout_r <= 12'h03F;
			12'hCA2 : dout_r <= 12'h03F;
			12'hCA3 : dout_r <= 12'h040;
			12'hCA4 : dout_r <= 12'h041;
			12'hCA5 : dout_r <= 12'h042;
			12'hCA6 : dout_r <= 12'h043;
			12'hCA7 : dout_r <= 12'h043;
			12'hCA8 : dout_r <= 12'h044;
			12'hCA9 : dout_r <= 12'h045;
			12'hCAA : dout_r <= 12'h046;
			12'hCAB : dout_r <= 12'h047;
			12'hCAC : dout_r <= 12'h047;
			12'hCAD : dout_r <= 12'h048;
			12'hCAE : dout_r <= 12'h049;
			12'hCAF : dout_r <= 12'h04A;
			12'hCB0 : dout_r <= 12'h04B;
			12'hCB1 : dout_r <= 12'h04B;
			12'hCB2 : dout_r <= 12'h04C;
			12'hCB3 : dout_r <= 12'h04D;
			12'hCB4 : dout_r <= 12'h04E;
			12'hCB5 : dout_r <= 12'h04F;
			12'hCB6 : dout_r <= 12'h050;
			12'hCB7 : dout_r <= 12'h051;
			12'hCB8 : dout_r <= 12'h051;
			12'hCB9 : dout_r <= 12'h052;
			12'hCBA : dout_r <= 12'h053;
			12'hCBB : dout_r <= 12'h054;
			12'hCBC : dout_r <= 12'h055;
			12'hCBD : dout_r <= 12'h056;
			12'hCBE : dout_r <= 12'h057;
			12'hCBF : dout_r <= 12'h058;
			12'hCC0 : dout_r <= 12'h059;
			12'hCC1 : dout_r <= 12'h05A;
			12'hCC2 : dout_r <= 12'h05A;
			12'hCC3 : dout_r <= 12'h05B;
			12'hCC4 : dout_r <= 12'h05C;
			12'hCC5 : dout_r <= 12'h05D;
			12'hCC6 : dout_r <= 12'h05E;
			12'hCC7 : dout_r <= 12'h05F;
			12'hCC8 : dout_r <= 12'h060;
			12'hCC9 : dout_r <= 12'h061;
			12'hCCA : dout_r <= 12'h062;
			12'hCCB : dout_r <= 12'h063;
			12'hCCC : dout_r <= 12'h064;
			12'hCCD : dout_r <= 12'h065;
			12'hCCE : dout_r <= 12'h066;
			12'hCCF : dout_r <= 12'h067;
			12'hCD0 : dout_r <= 12'h068;
			12'hCD1 : dout_r <= 12'h069;
			12'hCD2 : dout_r <= 12'h06A;
			12'hCD3 : dout_r <= 12'h06B;
			12'hCD4 : dout_r <= 12'h06C;
			12'hCD5 : dout_r <= 12'h06D;
			12'hCD6 : dout_r <= 12'h06E;
			12'hCD7 : dout_r <= 12'h06F;
			12'hCD8 : dout_r <= 12'h070;
			12'hCD9 : dout_r <= 12'h071;
			12'hCDA : dout_r <= 12'h072;
			12'hCDB : dout_r <= 12'h073;
			12'hCDC : dout_r <= 12'h074;
			12'hCDD : dout_r <= 12'h075;
			12'hCDE : dout_r <= 12'h076;
			12'hCDF : dout_r <= 12'h077;
			12'hCE0 : dout_r <= 12'h078;
			12'hCE1 : dout_r <= 12'h079;
			12'hCE2 : dout_r <= 12'h07A;
			12'hCE3 : dout_r <= 12'h07B;
			12'hCE4 : dout_r <= 12'h07C;
			12'hCE5 : dout_r <= 12'h07E;
			12'hCE6 : dout_r <= 12'h07F;
			12'hCE7 : dout_r <= 12'h080;
			12'hCE8 : dout_r <= 12'h081;
			12'hCE9 : dout_r <= 12'h082;
			12'hCEA : dout_r <= 12'h083;
			12'hCEB : dout_r <= 12'h084;
			12'hCEC : dout_r <= 12'h085;
			12'hCED : dout_r <= 12'h086;
			12'hCEE : dout_r <= 12'h087;
			12'hCEF : dout_r <= 12'h089;
			12'hCF0 : dout_r <= 12'h08A;
			12'hCF1 : dout_r <= 12'h08B;
			12'hCF2 : dout_r <= 12'h08C;
			12'hCF3 : dout_r <= 12'h08D;
			12'hCF4 : dout_r <= 12'h08E;
			12'hCF5 : dout_r <= 12'h08F;
			12'hCF6 : dout_r <= 12'h091;
			12'hCF7 : dout_r <= 12'h092;
			12'hCF8 : dout_r <= 12'h093;
			12'hCF9 : dout_r <= 12'h094;
			12'hCFA : dout_r <= 12'h095;
			12'hCFB : dout_r <= 12'h096;
			12'hCFC : dout_r <= 12'h098;
			12'hCFD : dout_r <= 12'h099;
			12'hCFE : dout_r <= 12'h09A;
			12'hCFF : dout_r <= 12'h09B;
			12'hD00 : dout_r <= 12'h09C;
			12'hD01 : dout_r <= 12'h09E;
			12'hD02 : dout_r <= 12'h09F;
			12'hD03 : dout_r <= 12'h0A0;
			12'hD04 : dout_r <= 12'h0A1;
			12'hD05 : dout_r <= 12'h0A2;
			12'hD06 : dout_r <= 12'h0A4;
			12'hD07 : dout_r <= 12'h0A5;
			12'hD08 : dout_r <= 12'h0A6;
			12'hD09 : dout_r <= 12'h0A7;
			12'hD0A : dout_r <= 12'h0A9;
			12'hD0B : dout_r <= 12'h0AA;
			12'hD0C : dout_r <= 12'h0AB;
			12'hD0D : dout_r <= 12'h0AC;
			12'hD0E : dout_r <= 12'h0AE;
			12'hD0F : dout_r <= 12'h0AF;
			12'hD10 : dout_r <= 12'h0B0;
			12'hD11 : dout_r <= 12'h0B1;
			12'hD12 : dout_r <= 12'h0B3;
			12'hD13 : dout_r <= 12'h0B4;
			12'hD14 : dout_r <= 12'h0B5;
			12'hD15 : dout_r <= 12'h0B7;
			12'hD16 : dout_r <= 12'h0B8;
			12'hD17 : dout_r <= 12'h0B9;
			12'hD18 : dout_r <= 12'h0BA;
			12'hD19 : dout_r <= 12'h0BC;
			12'hD1A : dout_r <= 12'h0BD;
			12'hD1B : dout_r <= 12'h0BE;
			12'hD1C : dout_r <= 12'h0C0;
			12'hD1D : dout_r <= 12'h0C1;
			12'hD1E : dout_r <= 12'h0C2;
			12'hD1F : dout_r <= 12'h0C4;
			12'hD20 : dout_r <= 12'h0C5;
			12'hD21 : dout_r <= 12'h0C6;
			12'hD22 : dout_r <= 12'h0C8;
			12'hD23 : dout_r <= 12'h0C9;
			12'hD24 : dout_r <= 12'h0CA;
			12'hD25 : dout_r <= 12'h0CC;
			12'hD26 : dout_r <= 12'h0CD;
			12'hD27 : dout_r <= 12'h0CF;
			12'hD28 : dout_r <= 12'h0D0;
			12'hD29 : dout_r <= 12'h0D1;
			12'hD2A : dout_r <= 12'h0D3;
			12'hD2B : dout_r <= 12'h0D4;
			12'hD2C : dout_r <= 12'h0D5;
			12'hD2D : dout_r <= 12'h0D7;
			12'hD2E : dout_r <= 12'h0D8;
			12'hD2F : dout_r <= 12'h0DA;
			12'hD30 : dout_r <= 12'h0DB;
			12'hD31 : dout_r <= 12'h0DC;
			12'hD32 : dout_r <= 12'h0DE;
			12'hD33 : dout_r <= 12'h0DF;
			12'hD34 : dout_r <= 12'h0E1;
			12'hD35 : dout_r <= 12'h0E2;
			12'hD36 : dout_r <= 12'h0E4;
			12'hD37 : dout_r <= 12'h0E5;
			12'hD38 : dout_r <= 12'h0E7;
			12'hD39 : dout_r <= 12'h0E8;
			12'hD3A : dout_r <= 12'h0E9;
			12'hD3B : dout_r <= 12'h0EB;
			12'hD3C : dout_r <= 12'h0EC;
			12'hD3D : dout_r <= 12'h0EE;
			12'hD3E : dout_r <= 12'h0EF;
			12'hD3F : dout_r <= 12'h0F1;
			12'hD40 : dout_r <= 12'h0F2;
			12'hD41 : dout_r <= 12'h0F4;
			12'hD42 : dout_r <= 12'h0F5;
			12'hD43 : dout_r <= 12'h0F7;
			12'hD44 : dout_r <= 12'h0F8;
			12'hD45 : dout_r <= 12'h0FA;
			12'hD46 : dout_r <= 12'h0FB;
			12'hD47 : dout_r <= 12'h0FD;
			12'hD48 : dout_r <= 12'h0FE;
			12'hD49 : dout_r <= 12'h100;
			12'hD4A : dout_r <= 12'h101;
			12'hD4B : dout_r <= 12'h103;
			12'hD4C : dout_r <= 12'h104;
			12'hD4D : dout_r <= 12'h106;
			12'hD4E : dout_r <= 12'h107;
			12'hD4F : dout_r <= 12'h109;
			12'hD50 : dout_r <= 12'h10A;
			12'hD51 : dout_r <= 12'h10C;
			12'hD52 : dout_r <= 12'h10E;
			12'hD53 : dout_r <= 12'h10F;
			12'hD54 : dout_r <= 12'h111;
			12'hD55 : dout_r <= 12'h112;
			12'hD56 : dout_r <= 12'h114;
			12'hD57 : dout_r <= 12'h115;
			12'hD58 : dout_r <= 12'h117;
			12'hD59 : dout_r <= 12'h119;
			12'hD5A : dout_r <= 12'h11A;
			12'hD5B : dout_r <= 12'h11C;
			12'hD5C : dout_r <= 12'h11D;
			12'hD5D : dout_r <= 12'h11F;
			12'hD5E : dout_r <= 12'h121;
			12'hD5F : dout_r <= 12'h122;
			12'hD60 : dout_r <= 12'h124;
			12'hD61 : dout_r <= 12'h125;
			12'hD62 : dout_r <= 12'h127;
			12'hD63 : dout_r <= 12'h129;
			12'hD64 : dout_r <= 12'h12A;
			12'hD65 : dout_r <= 12'h12C;
			12'hD66 : dout_r <= 12'h12D;
			12'hD67 : dout_r <= 12'h12F;
			12'hD68 : dout_r <= 12'h131;
			12'hD69 : dout_r <= 12'h132;
			12'hD6A : dout_r <= 12'h134;
			12'hD6B : dout_r <= 12'h136;
			12'hD6C : dout_r <= 12'h137;
			12'hD6D : dout_r <= 12'h139;
			12'hD6E : dout_r <= 12'h13B;
			12'hD6F : dout_r <= 12'h13C;
			12'hD70 : dout_r <= 12'h13E;
			12'hD71 : dout_r <= 12'h140;
			12'hD72 : dout_r <= 12'h141;
			12'hD73 : dout_r <= 12'h143;
			12'hD74 : dout_r <= 12'h145;
			12'hD75 : dout_r <= 12'h147;
			12'hD76 : dout_r <= 12'h148;
			12'hD77 : dout_r <= 12'h14A;
			12'hD78 : dout_r <= 12'h14C;
			12'hD79 : dout_r <= 12'h14D;
			12'hD7A : dout_r <= 12'h14F;
			12'hD7B : dout_r <= 12'h151;
			12'hD7C : dout_r <= 12'h153;
			12'hD7D : dout_r <= 12'h154;
			12'hD7E : dout_r <= 12'h156;
			12'hD7F : dout_r <= 12'h158;
			12'hD80 : dout_r <= 12'h159;
			12'hD81 : dout_r <= 12'h15B;
			12'hD82 : dout_r <= 12'h15D;
			12'hD83 : dout_r <= 12'h15F;
			12'hD84 : dout_r <= 12'h160;
			12'hD85 : dout_r <= 12'h162;
			12'hD86 : dout_r <= 12'h164;
			12'hD87 : dout_r <= 12'h166;
			12'hD88 : dout_r <= 12'h168;
			12'hD89 : dout_r <= 12'h169;
			12'hD8A : dout_r <= 12'h16B;
			12'hD8B : dout_r <= 12'h16D;
			12'hD8C : dout_r <= 12'h16F;
			12'hD8D : dout_r <= 12'h170;
			12'hD8E : dout_r <= 12'h172;
			12'hD8F : dout_r <= 12'h174;
			12'hD90 : dout_r <= 12'h176;
			12'hD91 : dout_r <= 12'h178;
			12'hD92 : dout_r <= 12'h17A;
			12'hD93 : dout_r <= 12'h17B;
			12'hD94 : dout_r <= 12'h17D;
			12'hD95 : dout_r <= 12'h17F;
			12'hD96 : dout_r <= 12'h181;
			12'hD97 : dout_r <= 12'h183;
			12'hD98 : dout_r <= 12'h184;
			12'hD99 : dout_r <= 12'h186;
			12'hD9A : dout_r <= 12'h188;
			12'hD9B : dout_r <= 12'h18A;
			12'hD9C : dout_r <= 12'h18C;
			12'hD9D : dout_r <= 12'h18E;
			12'hD9E : dout_r <= 12'h190;
			12'hD9F : dout_r <= 12'h191;
			12'hDA0 : dout_r <= 12'h193;
			12'hDA1 : dout_r <= 12'h195;
			12'hDA2 : dout_r <= 12'h197;
			12'hDA3 : dout_r <= 12'h199;
			12'hDA4 : dout_r <= 12'h19B;
			12'hDA5 : dout_r <= 12'h19D;
			12'hDA6 : dout_r <= 12'h19F;
			12'hDA7 : dout_r <= 12'h1A1;
			12'hDA8 : dout_r <= 12'h1A2;
			12'hDA9 : dout_r <= 12'h1A4;
			12'hDAA : dout_r <= 12'h1A6;
			12'hDAB : dout_r <= 12'h1A8;
			12'hDAC : dout_r <= 12'h1AA;
			12'hDAD : dout_r <= 12'h1AC;
			12'hDAE : dout_r <= 12'h1AE;
			12'hDAF : dout_r <= 12'h1B0;
			12'hDB0 : dout_r <= 12'h1B2;
			12'hDB1 : dout_r <= 12'h1B4;
			12'hDB2 : dout_r <= 12'h1B6;
			12'hDB3 : dout_r <= 12'h1B8;
			12'hDB4 : dout_r <= 12'h1BA;
			12'hDB5 : dout_r <= 12'h1BB;
			12'hDB6 : dout_r <= 12'h1BD;
			12'hDB7 : dout_r <= 12'h1BF;
			12'hDB8 : dout_r <= 12'h1C1;
			12'hDB9 : dout_r <= 12'h1C3;
			12'hDBA : dout_r <= 12'h1C5;
			12'hDBB : dout_r <= 12'h1C7;
			12'hDBC : dout_r <= 12'h1C9;
			12'hDBD : dout_r <= 12'h1CB;
			12'hDBE : dout_r <= 12'h1CD;
			12'hDBF : dout_r <= 12'h1CF;
			12'hDC0 : dout_r <= 12'h1D1;
			12'hDC1 : dout_r <= 12'h1D3;
			12'hDC2 : dout_r <= 12'h1D5;
			12'hDC3 : dout_r <= 12'h1D7;
			12'hDC4 : dout_r <= 12'h1D9;
			12'hDC5 : dout_r <= 12'h1DB;
			12'hDC6 : dout_r <= 12'h1DD;
			12'hDC7 : dout_r <= 12'h1DF;
			12'hDC8 : dout_r <= 12'h1E1;
			12'hDC9 : dout_r <= 12'h1E3;
			12'hDCA : dout_r <= 12'h1E5;
			12'hDCB : dout_r <= 12'h1E7;
			12'hDCC : dout_r <= 12'h1E9;
			12'hDCD : dout_r <= 12'h1EB;
			12'hDCE : dout_r <= 12'h1ED;
			12'hDCF : dout_r <= 12'h1EF;
			12'hDD0 : dout_r <= 12'h1F1;
			12'hDD1 : dout_r <= 12'h1F4;
			12'hDD2 : dout_r <= 12'h1F6;
			12'hDD3 : dout_r <= 12'h1F8;
			12'hDD4 : dout_r <= 12'h1FA;
			12'hDD5 : dout_r <= 12'h1FC;
			12'hDD6 : dout_r <= 12'h1FE;
			12'hDD7 : dout_r <= 12'h200;
			12'hDD8 : dout_r <= 12'h202;
			12'hDD9 : dout_r <= 12'h204;
			12'hDDA : dout_r <= 12'h206;
			12'hDDB : dout_r <= 12'h208;
			12'hDDC : dout_r <= 12'h20A;
			12'hDDD : dout_r <= 12'h20C;
			12'hDDE : dout_r <= 12'h20F;
			12'hDDF : dout_r <= 12'h211;
			12'hDE0 : dout_r <= 12'h213;
			12'hDE1 : dout_r <= 12'h215;
			12'hDE2 : dout_r <= 12'h217;
			12'hDE3 : dout_r <= 12'h219;
			12'hDE4 : dout_r <= 12'h21B;
			12'hDE5 : dout_r <= 12'h21D;
			12'hDE6 : dout_r <= 12'h21F;
			12'hDE7 : dout_r <= 12'h222;
			12'hDE8 : dout_r <= 12'h224;
			12'hDE9 : dout_r <= 12'h226;
			12'hDEA : dout_r <= 12'h228;
			12'hDEB : dout_r <= 12'h22A;
			12'hDEC : dout_r <= 12'h22C;
			12'hDED : dout_r <= 12'h22E;
			12'hDEE : dout_r <= 12'h231;
			12'hDEF : dout_r <= 12'h233;
			12'hDF0 : dout_r <= 12'h235;
			12'hDF1 : dout_r <= 12'h237;
			12'hDF2 : dout_r <= 12'h239;
			12'hDF3 : dout_r <= 12'h23B;
			12'hDF4 : dout_r <= 12'h23E;
			12'hDF5 : dout_r <= 12'h240;
			12'hDF6 : dout_r <= 12'h242;
			12'hDF7 : dout_r <= 12'h244;
			12'hDF8 : dout_r <= 12'h246;
			12'hDF9 : dout_r <= 12'h249;
			12'hDFA : dout_r <= 12'h24B;
			12'hDFB : dout_r <= 12'h24D;
			12'hDFC : dout_r <= 12'h24F;
			12'hDFD : dout_r <= 12'h251;
			12'hDFE : dout_r <= 12'h254;
			12'hDFF : dout_r <= 12'h256;
			12'hE00 : dout_r <= 12'h258;
			12'hE01 : dout_r <= 12'h25A;
			12'hE02 : dout_r <= 12'h25C;
			12'hE03 : dout_r <= 12'h25F;
			12'hE04 : dout_r <= 12'h261;
			12'hE05 : dout_r <= 12'h263;
			12'hE06 : dout_r <= 12'h265;
			12'hE07 : dout_r <= 12'h268;
			12'hE08 : dout_r <= 12'h26A;
			12'hE09 : dout_r <= 12'h26C;
			12'hE0A : dout_r <= 12'h26E;
			12'hE0B : dout_r <= 12'h271;
			12'hE0C : dout_r <= 12'h273;
			12'hE0D : dout_r <= 12'h275;
			12'hE0E : dout_r <= 12'h277;
			12'hE0F : dout_r <= 12'h27A;
			12'hE10 : dout_r <= 12'h27C;
			12'hE11 : dout_r <= 12'h27E;
			12'hE12 : dout_r <= 12'h281;
			12'hE13 : dout_r <= 12'h283;
			12'hE14 : dout_r <= 12'h285;
			12'hE15 : dout_r <= 12'h287;
			12'hE16 : dout_r <= 12'h28A;
			12'hE17 : dout_r <= 12'h28C;
			12'hE18 : dout_r <= 12'h28E;
			12'hE19 : dout_r <= 12'h291;
			12'hE1A : dout_r <= 12'h293;
			12'hE1B : dout_r <= 12'h295;
			12'hE1C : dout_r <= 12'h298;
			12'hE1D : dout_r <= 12'h29A;
			12'hE1E : dout_r <= 12'h29C;
			12'hE1F : dout_r <= 12'h29E;
			12'hE20 : dout_r <= 12'h2A1;
			12'hE21 : dout_r <= 12'h2A3;
			12'hE22 : dout_r <= 12'h2A5;
			12'hE23 : dout_r <= 12'h2A8;
			12'hE24 : dout_r <= 12'h2AA;
			12'hE25 : dout_r <= 12'h2AC;
			12'hE26 : dout_r <= 12'h2AF;
			12'hE27 : dout_r <= 12'h2B1;
			12'hE28 : dout_r <= 12'h2B4;
			12'hE29 : dout_r <= 12'h2B6;
			12'hE2A : dout_r <= 12'h2B8;
			12'hE2B : dout_r <= 12'h2BB;
			12'hE2C : dout_r <= 12'h2BD;
			12'hE2D : dout_r <= 12'h2BF;
			12'hE2E : dout_r <= 12'h2C2;
			12'hE2F : dout_r <= 12'h2C4;
			12'hE30 : dout_r <= 12'h2C6;
			12'hE31 : dout_r <= 12'h2C9;
			12'hE32 : dout_r <= 12'h2CB;
			12'hE33 : dout_r <= 12'h2CE;
			12'hE34 : dout_r <= 12'h2D0;
			12'hE35 : dout_r <= 12'h2D2;
			12'hE36 : dout_r <= 12'h2D5;
			12'hE37 : dout_r <= 12'h2D7;
			12'hE38 : dout_r <= 12'h2DA;
			12'hE39 : dout_r <= 12'h2DC;
			12'hE3A : dout_r <= 12'h2DE;
			12'hE3B : dout_r <= 12'h2E1;
			12'hE3C : dout_r <= 12'h2E3;
			12'hE3D : dout_r <= 12'h2E6;
			12'hE3E : dout_r <= 12'h2E8;
			12'hE3F : dout_r <= 12'h2EA;
			12'hE40 : dout_r <= 12'h2ED;
			12'hE41 : dout_r <= 12'h2EF;
			12'hE42 : dout_r <= 12'h2F2;
			12'hE43 : dout_r <= 12'h2F4;
			12'hE44 : dout_r <= 12'h2F7;
			12'hE45 : dout_r <= 12'h2F9;
			12'hE46 : dout_r <= 12'h2FC;
			12'hE47 : dout_r <= 12'h2FE;
			12'hE48 : dout_r <= 12'h300;
			12'hE49 : dout_r <= 12'h303;
			12'hE4A : dout_r <= 12'h305;
			12'hE4B : dout_r <= 12'h308;
			12'hE4C : dout_r <= 12'h30A;
			12'hE4D : dout_r <= 12'h30D;
			12'hE4E : dout_r <= 12'h30F;
			12'hE4F : dout_r <= 12'h312;
			12'hE50 : dout_r <= 12'h314;
			12'hE51 : dout_r <= 12'h317;
			12'hE52 : dout_r <= 12'h319;
			12'hE53 : dout_r <= 12'h31C;
			12'hE54 : dout_r <= 12'h31E;
			12'hE55 : dout_r <= 12'h321;
			12'hE56 : dout_r <= 12'h323;
			12'hE57 : dout_r <= 12'h326;
			12'hE58 : dout_r <= 12'h328;
			12'hE59 : dout_r <= 12'h32B;
			12'hE5A : dout_r <= 12'h32D;
			12'hE5B : dout_r <= 12'h330;
			12'hE5C : dout_r <= 12'h332;
			12'hE5D : dout_r <= 12'h335;
			12'hE5E : dout_r <= 12'h337;
			12'hE5F : dout_r <= 12'h33A;
			12'hE60 : dout_r <= 12'h33C;
			12'hE61 : dout_r <= 12'h33F;
			12'hE62 : dout_r <= 12'h341;
			12'hE63 : dout_r <= 12'h344;
			12'hE64 : dout_r <= 12'h346;
			12'hE65 : dout_r <= 12'h349;
			12'hE66 : dout_r <= 12'h34B;
			12'hE67 : dout_r <= 12'h34E;
			12'hE68 : dout_r <= 12'h350;
			12'hE69 : dout_r <= 12'h353;
			12'hE6A : dout_r <= 12'h355;
			12'hE6B : dout_r <= 12'h358;
			12'hE6C : dout_r <= 12'h35B;
			12'hE6D : dout_r <= 12'h35D;
			12'hE6E : dout_r <= 12'h360;
			12'hE6F : dout_r <= 12'h362;
			12'hE70 : dout_r <= 12'h365;
			12'hE71 : dout_r <= 12'h367;
			12'hE72 : dout_r <= 12'h36A;
			12'hE73 : dout_r <= 12'h36D;
			12'hE74 : dout_r <= 12'h36F;
			12'hE75 : dout_r <= 12'h372;
			12'hE76 : dout_r <= 12'h374;
			12'hE77 : dout_r <= 12'h377;
			12'hE78 : dout_r <= 12'h379;
			12'hE79 : dout_r <= 12'h37C;
			12'hE7A : dout_r <= 12'h37F;
			12'hE7B : dout_r <= 12'h381;
			12'hE7C : dout_r <= 12'h384;
			12'hE7D : dout_r <= 12'h386;
			12'hE7E : dout_r <= 12'h389;
			12'hE7F : dout_r <= 12'h38C;
			12'hE80 : dout_r <= 12'h38E;
			12'hE81 : dout_r <= 12'h391;
			12'hE82 : dout_r <= 12'h393;
			12'hE83 : dout_r <= 12'h396;
			12'hE84 : dout_r <= 12'h399;
			12'hE85 : dout_r <= 12'h39B;
			12'hE86 : dout_r <= 12'h39E;
			12'hE87 : dout_r <= 12'h3A1;
			12'hE88 : dout_r <= 12'h3A3;
			12'hE89 : dout_r <= 12'h3A6;
			12'hE8A : dout_r <= 12'h3A8;
			12'hE8B : dout_r <= 12'h3AB;
			12'hE8C : dout_r <= 12'h3AE;
			12'hE8D : dout_r <= 12'h3B0;
			12'hE8E : dout_r <= 12'h3B3;
			12'hE8F : dout_r <= 12'h3B6;
			12'hE90 : dout_r <= 12'h3B8;
			12'hE91 : dout_r <= 12'h3BB;
			12'hE92 : dout_r <= 12'h3BE;
			12'hE93 : dout_r <= 12'h3C0;
			12'hE94 : dout_r <= 12'h3C3;
			12'hE95 : dout_r <= 12'h3C6;
			12'hE96 : dout_r <= 12'h3C8;
			12'hE97 : dout_r <= 12'h3CB;
			12'hE98 : dout_r <= 12'h3CE;
			12'hE99 : dout_r <= 12'h3D0;
			12'hE9A : dout_r <= 12'h3D3;
			12'hE9B : dout_r <= 12'h3D6;
			12'hE9C : dout_r <= 12'h3D8;
			12'hE9D : dout_r <= 12'h3DB;
			12'hE9E : dout_r <= 12'h3DE;
			12'hE9F : dout_r <= 12'h3E0;
			12'hEA0 : dout_r <= 12'h3E3;
			12'hEA1 : dout_r <= 12'h3E6;
			12'hEA2 : dout_r <= 12'h3E9;
			12'hEA3 : dout_r <= 12'h3EB;
			12'hEA4 : dout_r <= 12'h3EE;
			12'hEA5 : dout_r <= 12'h3F1;
			12'hEA6 : dout_r <= 12'h3F3;
			12'hEA7 : dout_r <= 12'h3F6;
			12'hEA8 : dout_r <= 12'h3F9;
			12'hEA9 : dout_r <= 12'h3FB;
			12'hEAA : dout_r <= 12'h3FE;
			12'hEAB : dout_r <= 12'h401;
			12'hEAC : dout_r <= 12'h404;
			12'hEAD : dout_r <= 12'h406;
			12'hEAE : dout_r <= 12'h409;
			12'hEAF : dout_r <= 12'h40C;
			12'hEB0 : dout_r <= 12'h40F;
			12'hEB1 : dout_r <= 12'h411;
			12'hEB2 : dout_r <= 12'h414;
			12'hEB3 : dout_r <= 12'h417;
			12'hEB4 : dout_r <= 12'h419;
			12'hEB5 : dout_r <= 12'h41C;
			12'hEB6 : dout_r <= 12'h41F;
			12'hEB7 : dout_r <= 12'h422;
			12'hEB8 : dout_r <= 12'h424;
			12'hEB9 : dout_r <= 12'h427;
			12'hEBA : dout_r <= 12'h42A;
			12'hEBB : dout_r <= 12'h42D;
			12'hEBC : dout_r <= 12'h42F;
			12'hEBD : dout_r <= 12'h432;
			12'hEBE : dout_r <= 12'h435;
			12'hEBF : dout_r <= 12'h438;
			12'hEC0 : dout_r <= 12'h43B;
			12'hEC1 : dout_r <= 12'h43D;
			12'hEC2 : dout_r <= 12'h440;
			12'hEC3 : dout_r <= 12'h443;
			12'hEC4 : dout_r <= 12'h446;
			12'hEC5 : dout_r <= 12'h448;
			12'hEC6 : dout_r <= 12'h44B;
			12'hEC7 : dout_r <= 12'h44E;
			12'hEC8 : dout_r <= 12'h451;
			12'hEC9 : dout_r <= 12'h454;
			12'hECA : dout_r <= 12'h456;
			12'hECB : dout_r <= 12'h459;
			12'hECC : dout_r <= 12'h45C;
			12'hECD : dout_r <= 12'h45F;
			12'hECE : dout_r <= 12'h462;
			12'hECF : dout_r <= 12'h464;
			12'hED0 : dout_r <= 12'h467;
			12'hED1 : dout_r <= 12'h46A;
			12'hED2 : dout_r <= 12'h46D;
			12'hED3 : dout_r <= 12'h470;
			12'hED4 : dout_r <= 12'h472;
			12'hED5 : dout_r <= 12'h475;
			12'hED6 : dout_r <= 12'h478;
			12'hED7 : dout_r <= 12'h47B;
			12'hED8 : dout_r <= 12'h47E;
			12'hED9 : dout_r <= 12'h480;
			12'hEDA : dout_r <= 12'h483;
			12'hEDB : dout_r <= 12'h486;
			12'hEDC : dout_r <= 12'h489;
			12'hEDD : dout_r <= 12'h48C;
			12'hEDE : dout_r <= 12'h48F;
			12'hEDF : dout_r <= 12'h491;
			12'hEE0 : dout_r <= 12'h494;
			12'hEE1 : dout_r <= 12'h497;
			12'hEE2 : dout_r <= 12'h49A;
			12'hEE3 : dout_r <= 12'h49D;
			12'hEE4 : dout_r <= 12'h4A0;
			12'hEE5 : dout_r <= 12'h4A3;
			12'hEE6 : dout_r <= 12'h4A5;
			12'hEE7 : dout_r <= 12'h4A8;
			12'hEE8 : dout_r <= 12'h4AB;
			12'hEE9 : dout_r <= 12'h4AE;
			12'hEEA : dout_r <= 12'h4B1;
			12'hEEB : dout_r <= 12'h4B4;
			12'hEEC : dout_r <= 12'h4B7;
			12'hEED : dout_r <= 12'h4B9;
			12'hEEE : dout_r <= 12'h4BC;
			12'hEEF : dout_r <= 12'h4BF;
			12'hEF0 : dout_r <= 12'h4C2;
			12'hEF1 : dout_r <= 12'h4C5;
			12'hEF2 : dout_r <= 12'h4C8;
			12'hEF3 : dout_r <= 12'h4CB;
			12'hEF4 : dout_r <= 12'h4CD;
			12'hEF5 : dout_r <= 12'h4D0;
			12'hEF6 : dout_r <= 12'h4D3;
			12'hEF7 : dout_r <= 12'h4D6;
			12'hEF8 : dout_r <= 12'h4D9;
			12'hEF9 : dout_r <= 12'h4DC;
			12'hEFA : dout_r <= 12'h4DF;
			12'hEFB : dout_r <= 12'h4E2;
			12'hEFC : dout_r <= 12'h4E5;
			12'hEFD : dout_r <= 12'h4E7;
			12'hEFE : dout_r <= 12'h4EA;
			12'hEFF : dout_r <= 12'h4ED;
			12'hF00 : dout_r <= 12'h4F0;
			12'hF01 : dout_r <= 12'h4F3;
			12'hF02 : dout_r <= 12'h4F6;
			12'hF03 : dout_r <= 12'h4F9;
			12'hF04 : dout_r <= 12'h4FC;
			12'hF05 : dout_r <= 12'h4FF;
			12'hF06 : dout_r <= 12'h502;
			12'hF07 : dout_r <= 12'h504;
			12'hF08 : dout_r <= 12'h507;
			12'hF09 : dout_r <= 12'h50A;
			12'hF0A : dout_r <= 12'h50D;
			12'hF0B : dout_r <= 12'h510;
			12'hF0C : dout_r <= 12'h513;
			12'hF0D : dout_r <= 12'h516;
			12'hF0E : dout_r <= 12'h519;
			12'hF0F : dout_r <= 12'h51C;
			12'hF10 : dout_r <= 12'h51F;
			12'hF11 : dout_r <= 12'h522;
			12'hF12 : dout_r <= 12'h525;
			12'hF13 : dout_r <= 12'h528;
			12'hF14 : dout_r <= 12'h52B;
			12'hF15 : dout_r <= 12'h52D;
			12'hF16 : dout_r <= 12'h530;
			12'hF17 : dout_r <= 12'h533;
			12'hF18 : dout_r <= 12'h536;
			12'hF19 : dout_r <= 12'h539;
			12'hF1A : dout_r <= 12'h53C;
			12'hF1B : dout_r <= 12'h53F;
			12'hF1C : dout_r <= 12'h542;
			12'hF1D : dout_r <= 12'h545;
			12'hF1E : dout_r <= 12'h548;
			12'hF1F : dout_r <= 12'h54B;
			12'hF20 : dout_r <= 12'h54E;
			12'hF21 : dout_r <= 12'h551;
			12'hF22 : dout_r <= 12'h554;
			12'hF23 : dout_r <= 12'h557;
			12'hF24 : dout_r <= 12'h55A;
			12'hF25 : dout_r <= 12'h55D;
			12'hF26 : dout_r <= 12'h560;
			12'hF27 : dout_r <= 12'h563;
			12'hF28 : dout_r <= 12'h566;
			12'hF29 : dout_r <= 12'h569;
			12'hF2A : dout_r <= 12'h56C;
			12'hF2B : dout_r <= 12'h56F;
			12'hF2C : dout_r <= 12'h571;
			12'hF2D : dout_r <= 12'h574;
			12'hF2E : dout_r <= 12'h577;
			12'hF2F : dout_r <= 12'h57A;
			12'hF30 : dout_r <= 12'h57D;
			12'hF31 : dout_r <= 12'h580;
			12'hF32 : dout_r <= 12'h583;
			12'hF33 : dout_r <= 12'h586;
			12'hF34 : dout_r <= 12'h589;
			12'hF35 : dout_r <= 12'h58C;
			12'hF36 : dout_r <= 12'h58F;
			12'hF37 : dout_r <= 12'h592;
			12'hF38 : dout_r <= 12'h595;
			12'hF39 : dout_r <= 12'h598;
			12'hF3A : dout_r <= 12'h59B;
			12'hF3B : dout_r <= 12'h59E;
			12'hF3C : dout_r <= 12'h5A1;
			12'hF3D : dout_r <= 12'h5A4;
			12'hF3E : dout_r <= 12'h5A7;
			12'hF3F : dout_r <= 12'h5AA;
			12'hF40 : dout_r <= 12'h5AD;
			12'hF41 : dout_r <= 12'h5B0;
			12'hF42 : dout_r <= 12'h5B3;
			12'hF43 : dout_r <= 12'h5B6;
			12'hF44 : dout_r <= 12'h5B9;
			12'hF45 : dout_r <= 12'h5BC;
			12'hF46 : dout_r <= 12'h5BF;
			12'hF47 : dout_r <= 12'h5C2;
			12'hF48 : dout_r <= 12'h5C5;
			12'hF49 : dout_r <= 12'h5C8;
			12'hF4A : dout_r <= 12'h5CB;
			12'hF4B : dout_r <= 12'h5CE;
			12'hF4C : dout_r <= 12'h5D1;
			12'hF4D : dout_r <= 12'h5D4;
			12'hF4E : dout_r <= 12'h5D7;
			12'hF4F : dout_r <= 12'h5DB;
			12'hF50 : dout_r <= 12'h5DE;
			12'hF51 : dout_r <= 12'h5E1;
			12'hF52 : dout_r <= 12'h5E4;
			12'hF53 : dout_r <= 12'h5E7;
			12'hF54 : dout_r <= 12'h5EA;
			12'hF55 : dout_r <= 12'h5ED;
			12'hF56 : dout_r <= 12'h5F0;
			12'hF57 : dout_r <= 12'h5F3;
			12'hF58 : dout_r <= 12'h5F6;
			12'hF59 : dout_r <= 12'h5F9;
			12'hF5A : dout_r <= 12'h5FC;
			12'hF5B : dout_r <= 12'h5FF;
			12'hF5C : dout_r <= 12'h602;
			12'hF5D : dout_r <= 12'h605;
			12'hF5E : dout_r <= 12'h608;
			12'hF5F : dout_r <= 12'h60B;
			12'hF60 : dout_r <= 12'h60E;
			12'hF61 : dout_r <= 12'h611;
			12'hF62 : dout_r <= 12'h614;
			12'hF63 : dout_r <= 12'h617;
			12'hF64 : dout_r <= 12'h61A;
			12'hF65 : dout_r <= 12'h61D;
			12'hF66 : dout_r <= 12'h620;
			12'hF67 : dout_r <= 12'h623;
			12'hF68 : dout_r <= 12'h627;
			12'hF69 : dout_r <= 12'h62A;
			12'hF6A : dout_r <= 12'h62D;
			12'hF6B : dout_r <= 12'h630;
			12'hF6C : dout_r <= 12'h633;
			12'hF6D : dout_r <= 12'h636;
			12'hF6E : dout_r <= 12'h639;
			12'hF6F : dout_r <= 12'h63C;
			12'hF70 : dout_r <= 12'h63F;
			12'hF71 : dout_r <= 12'h642;
			12'hF72 : dout_r <= 12'h645;
			12'hF73 : dout_r <= 12'h648;
			12'hF74 : dout_r <= 12'h64B;
			12'hF75 : dout_r <= 12'h64E;
			12'hF76 : dout_r <= 12'h651;
			12'hF77 : dout_r <= 12'h654;
			12'hF78 : dout_r <= 12'h658;
			12'hF79 : dout_r <= 12'h65B;
			12'hF7A : dout_r <= 12'h65E;
			12'hF7B : dout_r <= 12'h661;
			12'hF7C : dout_r <= 12'h664;
			12'hF7D : dout_r <= 12'h667;
			12'hF7E : dout_r <= 12'h66A;
			12'hF7F : dout_r <= 12'h66D;
			12'hF80 : dout_r <= 12'h670;
			12'hF81 : dout_r <= 12'h673;
			12'hF82 : dout_r <= 12'h676;
			12'hF83 : dout_r <= 12'h679;
			12'hF84 : dout_r <= 12'h67C;
			12'hF85 : dout_r <= 12'h680;
			12'hF86 : dout_r <= 12'h683;
			12'hF87 : dout_r <= 12'h686;
			12'hF88 : dout_r <= 12'h689;
			12'hF89 : dout_r <= 12'h68C;
			12'hF8A : dout_r <= 12'h68F;
			12'hF8B : dout_r <= 12'h692;
			12'hF8C : dout_r <= 12'h695;
			12'hF8D : dout_r <= 12'h698;
			12'hF8E : dout_r <= 12'h69B;
			12'hF8F : dout_r <= 12'h69E;
			12'hF90 : dout_r <= 12'h6A2;
			12'hF91 : dout_r <= 12'h6A5;
			12'hF92 : dout_r <= 12'h6A8;
			12'hF93 : dout_r <= 12'h6AB;
			12'hF94 : dout_r <= 12'h6AE;
			12'hF95 : dout_r <= 12'h6B1;
			12'hF96 : dout_r <= 12'h6B4;
			12'hF97 : dout_r <= 12'h6B7;
			12'hF98 : dout_r <= 12'h6BA;
			12'hF99 : dout_r <= 12'h6BD;
			12'hF9A : dout_r <= 12'h6C1;
			12'hF9B : dout_r <= 12'h6C4;
			12'hF9C : dout_r <= 12'h6C7;
			12'hF9D : dout_r <= 12'h6CA;
			12'hF9E : dout_r <= 12'h6CD;
			12'hF9F : dout_r <= 12'h6D0;
			12'hFA0 : dout_r <= 12'h6D3;
			12'hFA1 : dout_r <= 12'h6D6;
			12'hFA2 : dout_r <= 12'h6D9;
			12'hFA3 : dout_r <= 12'h6DC;
			12'hFA4 : dout_r <= 12'h6E0;
			12'hFA5 : dout_r <= 12'h6E3;
			12'hFA6 : dout_r <= 12'h6E6;
			12'hFA7 : dout_r <= 12'h6E9;
			12'hFA8 : dout_r <= 12'h6EC;
			12'hFA9 : dout_r <= 12'h6EF;
			12'hFAA : dout_r <= 12'h6F2;
			12'hFAB : dout_r <= 12'h6F5;
			12'hFAC : dout_r <= 12'h6F8;
			12'hFAD : dout_r <= 12'h6FC;
			12'hFAE : dout_r <= 12'h6FF;
			12'hFAF : dout_r <= 12'h702;
			12'hFB0 : dout_r <= 12'h705;
			12'hFB1 : dout_r <= 12'h708;
			12'hFB2 : dout_r <= 12'h70B;
			12'hFB3 : dout_r <= 12'h70E;
			12'hFB4 : dout_r <= 12'h711;
			12'hFB5 : dout_r <= 12'h715;
			12'hFB6 : dout_r <= 12'h718;
			12'hFB7 : dout_r <= 12'h71B;
			12'hFB8 : dout_r <= 12'h71E;
			12'hFB9 : dout_r <= 12'h721;
			12'hFBA : dout_r <= 12'h724;
			12'hFBB : dout_r <= 12'h727;
			12'hFBC : dout_r <= 12'h72A;
			12'hFBD : dout_r <= 12'h72D;
			12'hFBE : dout_r <= 12'h731;
			12'hFBF : dout_r <= 12'h734;
			12'hFC0 : dout_r <= 12'h737;
			12'hFC1 : dout_r <= 12'h73A;
			12'hFC2 : dout_r <= 12'h73D;
			12'hFC3 : dout_r <= 12'h740;
			12'hFC4 : dout_r <= 12'h743;
			12'hFC5 : dout_r <= 12'h746;
			12'hFC6 : dout_r <= 12'h74A;
			12'hFC7 : dout_r <= 12'h74D;
			12'hFC8 : dout_r <= 12'h750;
			12'hFC9 : dout_r <= 12'h753;
			12'hFCA : dout_r <= 12'h756;
			12'hFCB : dout_r <= 12'h759;
			12'hFCC : dout_r <= 12'h75C;
			12'hFCD : dout_r <= 12'h760;
			12'hFCE : dout_r <= 12'h763;
			12'hFCF : dout_r <= 12'h766;
			12'hFD0 : dout_r <= 12'h769;
			12'hFD1 : dout_r <= 12'h76C;
			12'hFD2 : dout_r <= 12'h76F;
			12'hFD3 : dout_r <= 12'h772;
			12'hFD4 : dout_r <= 12'h775;
			12'hFD5 : dout_r <= 12'h779;
			12'hFD6 : dout_r <= 12'h77C;
			12'hFD7 : dout_r <= 12'h77F;
			12'hFD8 : dout_r <= 12'h782;
			12'hFD9 : dout_r <= 12'h785;
			12'hFDA : dout_r <= 12'h788;
			12'hFDB : dout_r <= 12'h78B;
			12'hFDC : dout_r <= 12'h78F;
			12'hFDD : dout_r <= 12'h792;
			12'hFDE : dout_r <= 12'h795;
			12'hFDF : dout_r <= 12'h798;
			12'hFE0 : dout_r <= 12'h79B;
			12'hFE1 : dout_r <= 12'h79E;
			12'hFE2 : dout_r <= 12'h7A1;
			12'hFE3 : dout_r <= 12'h7A4;
			12'hFE4 : dout_r <= 12'h7A8;
			12'hFE5 : dout_r <= 12'h7AB;
			12'hFE6 : dout_r <= 12'h7AE;
			12'hFE7 : dout_r <= 12'h7B1;
			12'hFE8 : dout_r <= 12'h7B4;
			12'hFE9 : dout_r <= 12'h7B7;
			12'hFEA : dout_r <= 12'h7BA;
			12'hFEB : dout_r <= 12'h7BE;
			12'hFEC : dout_r <= 12'h7C1;
			12'hFED : dout_r <= 12'h7C4;
			12'hFEE : dout_r <= 12'h7C7;
			12'hFEF : dout_r <= 12'h7CA;
			12'hFF0 : dout_r <= 12'h7CD;
			12'hFF1 : dout_r <= 12'h7D0;
			12'hFF2 : dout_r <= 12'h7D4;
			12'hFF3 : dout_r <= 12'h7D7;
			12'hFF4 : dout_r <= 12'h7DA;
			12'hFF5 : dout_r <= 12'h7DD;
			12'hFF6 : dout_r <= 12'h7E0;
			12'hFF7 : dout_r <= 12'h7E3;
			12'hFF8 : dout_r <= 12'h7E6;
			12'hFF9 : dout_r <= 12'h7EA;
			12'hFFA : dout_r <= 12'h7ED;
			12'hFFB : dout_r <= 12'h7F0;
			12'hFFC : dout_r <= 12'h7F3;
			12'hFFD : dout_r <= 12'h7F6;
			12'hFFE : dout_r <= 12'h7F9;
			12'hFFF : dout_r <= 12'h7FC;
			endcase
	end	

	//wire output
	assign dout = dout_r;
	
endmodule
